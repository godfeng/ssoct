��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� (� ��"fف�����͎��T�k ������[���a�8%`��4�s�6�XAoeu��a@����þ�V�\O����L�N��<G� �mD�?ea�8�����B}rs4��������b�N<��;��� B]�pE���	x]̃Dj#^Da����M�ٲ��9ߪ�
�M��ļz����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω�[@�qR�� (� ��"fف�����͎��T�k ���������	x]̢/����w�c.$���S���bJ���<����PГ����"��N�� <9[�8@������G�٘���ty.hSN�����\�4�smg�:�TZz�0Q�����F���0FUR�.�;�~�MUs �P�^,�Q����j�_��l�؊9��8���M�3)ͰnL
�k�8���҆�|n������}�K-���W}��@_���J�Й�m����u�����w`q�tc�ؑ��g�=Iĩ�m��d�7�Q����.P2:}��>�,�_'�hQr�k@Q��j��C�뫰v]uR����Pl����N�Er��xXc)O�%���ʅ�$n��RL�a)�ƞ��U<���G�/9Ɗ���ބ�F=��?�r�7C��H���j�v�?��$m��2߼
�d�
 O4�J�|(�����	x]�<���eo�l$����Pfg��w{��������PГ��-�������n�GE^��.�Ū�'E���f!ۤՀ/Q9*سBK-����s~�j1���u��w)�S �J���vy�~篟|�<8�F�-:�0��E_}�8�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A`�6��{���9��m�!=�y����h�}�N�5�%��/��Hg2�5��o?�M��;]���>��G�0��H��k3��Ԩr�`����ǆjqcA�f�J��p�E��PN!y�(�����g�v-���I?���l����P=�����S��@�"G�C�(�%A��I�\��M���~'B>��B_���� Z�X�U�e0���0�vs�6��g.zQ��!K�4����\�4�s��{��]Qǯ�����ջ���­�WSt!K� �~�MUs H6).���o�6=� �wx0�<�����%���Z�G�a}C��aA�O�Yv������}�N�n��ՙ����
-�k�8���҆�|n����0ӵ*4�I�(ۿ�az|U�J�Й�m��\�e	���ȏ=���Y�*/�o)�>Ճ3��5�2G�$&��@�r�<ؔC95^T�,+Ⱦ
� �AH�����`�y$h��ݔf5*`]�mV�W���ڇ~�MUs c�+պNE��#Y��#p��'��������S�����:�֣I���Y/��S"�:����:�wl B����/��;��|B�6L����k�y.�)$����\�4�sm�|E ,mߍu�M9ts{z>�z�J�S��6CL�7C��H!�������0�"���L�M�=o����"���	x]�9ڿ��Qc�J�M=��t�R���:�ڣԏ�8�:r&@/_�x{�֐@����)���h=��&��C_�m�!=�y����h�}�G���AjD7Z����~�<�*h�u���;����K�@�c$�S�in���ћ�A����ȧг'?��j���}�?�����ל��*����	� D����	��\�4�slom��Qjh�6g��c���w�]� ܩ�*�o?�M��;]�NT[�=� ����i�D���_i��Z��71��%�}Ř&�� �W�#!��Y�:pRр��>�B�m�!=�y����h�}ۨ���'_I2���|����=T�k�u���;��o��&`o�3�P2��]�:��0��H��k3��ԨrZ��U��+@G�1����RL�a)�G{�<����I��V�Sn��t>�h�9!�zg�Z�$�%dZ&��Ǯ"�lf�~��m���w>�K�6���	x]�m�Je{q��N��(
{��DIU�J���<���&}Xa���������dG�b�{����V���	x]���Ec��$7��Mv�9��!��|�PS��N8�:r&@㽕����u�f�W��}ƪ%I/ο��굶m�!=�y����h�}jh�6g������\��>1�ij��o?�M��;]M�ֲ,�� �`���ё�?��9)I����C��
� �AH�)��H�� �b5z����;���8l�TS�F@�4%��%dZ&��Ǯ"�lf�~��m���w>�K�6���	x]̍��;������,b�S�����w{����֩��jR�"�H�ٳ,�M(F�N��d�>�l;��r�O��C��0��$�>��w�!�S�?|eU�����u���;��ü	A�3��<�ؒHXڏ`ϥK� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S)�-E����}����E���ƪ�(����D�I�?g�f� gt~��~)�-E��r���q P�^�&d�A|�1�:�Ω��
�/�r�ѬL�1m��+5z�P�_X�I�?g�f�$��P��� �}E+���c�W_QL�ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l�������+rb����Uh7u+��T��٤�2[51g~Ӝ��ajƎ�c��(r���U����+rb��{b�2"��-h|,���(����>S��ә�����/�4�}n'���a*�x���� ����ޙB!7����ˉ�1�:�Ω�[@�qR�� (� ��"fف�����Z�NCIw4t�iZ]XF�������� ��k\�\�KE���H���o��qo�:�ȓ��o)�]r k�|6�8��u*K6H.��h��u>j޽���Ǜ������[7�d|���XP��Ȩ�wl��h�Vx�%L��Ok��@zL͊�q���Vǃ���G&%	��ڔ��n����\�v�)��+�}��]�.�b�;װ?�p��U��֜��3JHn��z���G7�����o)�]rN�ǁ�f�T�J��H9��\�v�T?�7G|`^�R@Κ�2�Ix���KaJuA�����IÙ=�HF���m¡�3
�v�v-}�	mp�EN��S�IÙ=�H%v@����fnQ�rV4����X���\�v���GAџV^�R@Κ�2'�̗������\�ݠ�3zL͊�q��UG�s�����M���o�G�m�?M�*B�[zL͊�q��UG�s�����M���HaU$kX��� nU�IÙ=�HF���m¡A�h��+Fen����9��#�B�sYC��\�v��_�R�G�$����{v��G�K$xE�p4rqG7��u*K6H �i7�sp>��%��H��5[�����q�_�N�6�Ặ��Ϊ�Q� ~�����(��q�
�Bk�i�E?�xu����ma��u��ۯi\�q���Ì �&�k��>���c��d�|ݔ�3�5�}�]���x�]�V�����Ү��`�+S�p��ͷQ�X����fx'v�ao.\C�k�ף�D�~4#C(�}�IÙ=�H�%��@�Kǹ|���|u��RJHn��z��r9�3��X�u�ӑ�띂ii�4];ˍH���Vchw�D��y.���=��܄��띂ii�4];ˍH���Vchw�D��y.���eŞG�T(x�]�V���o��8���Cf֩Q�e]��W�'NTؕ@�.MŃ�,��)x�]�V���F�uB�W˪��/h�Б����x�]�V��,t����t�i�lK�I<��fҾ��9��ЂDa��(o��0��7��|g�Y�'���Xw�f�VHF��Q�#<4^�v�ј�"��Z鎬����F�71�B�������%�N�By3��<�]�!����M[��Ǣ�L ʞ��0��m��x���j���0z�cUL3�X�j��7$2Ӕ�1���_�wa(􆿳�tP"7��%e��0�U+�qbp@��wbk�$���7Z���(�
t�ژq���U� бb*	��|	�WI�����
L'���Xw�4��}�<�=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A����ɻ:�E�1N�By3��<�]�!���\B��V���#���L�
�����Yl���#�]�!��	Ǹ�y85��(�C)&���lC��U�T�\ �͹g}|�H���p��b��e������]�!��	Ǹ�y85���ǳ@�M�H�ɇM��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+�ڔ�wV��y�p�cP ������w�f�����67�a��c���}��D���(��z�j�)�q��1�:�Ω�[@�qR�� (� ��"fف�����Z�NCIw4C#/<���q�]��`4Ƹp�iF��6P�;ń�X�����64B�su� Z�O )�\�~xy�}w˙��2����1�~�+��E"!o���]	��Ptb(Sl�z=�y:D���';:ZËF�3$����Vܙ���LM �EVܕ����������a�"�'n�^0ohC$?���;���EWr��uNS\IÙ=�H1�Z8[iI9�o����"��y�S�yH��"J�A��S+B�l�^>*���a�"�_���3��q�l;1����bU�򍬓BS���Usdx����p��nk�R���c&;�L�FZ�1Ǩ�Yc�A�/����<.+6J!�5����`Kְ�4'N5wĒ����H���o��qo�:���$��Xo���~��1�51	�<�����ȳ�%�MZẶ��Ϊ���Jjz�p�m~|�֛� �>��h �=��b9����lY1�ËF�3$����Vܙ���n%�G�33p�m~|����� �ܰ�a\Y����+���LQ��b9������U.6��̞��>��3
�v�v-}�	mp@�s�p���.ᬵy���"�n��T̞��>�h�5,Wlr�r%)cA��gx�܈�5����`Kss2����`�|��K�z�!��(�����3xļ�\�v�o���H�|k��!a�tc�&ck�����1ٞ<h���/��&�[�$��X�>��u��>п�p=	�˳͠m�xW��9u$d9��}ϔ��J�s���
�k��!a�tc�&ck��°������R�wX�����/��&�[�$��X�S�wS& >ht[�����GI$��ǂcY�~�s<��MR�ɧ�	tc&�j��1�a-���7a
��r����~v����"X��[��Q[R�7��z�h��4�*ܑe�W����n�4�c_����+.�	|ǔ�.Yz�Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P�|h{�T��`�)�	�%{�;���;�L���9o��+hi�?O��K�����=ў@'���Xw�j�7��Vx�%L��W��_�ړ8���/��֍z����I��'�ct�:��RE�QS����>�b9���S�nU�&u������u��U|<��⏇���;�z*���Be�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�F�������T�\ �͠ �ݺ��I��'�������.��R�}vJ^�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xǩ"�4s2nQ�rV� �L_K�*��M���HaU$kX�GY�=�=T������.��R�}vJ^*h�!<^�5����`K݁.�q�0��E|�,1#��Z����_c��(���B��j�Q��9�V�ݦ\�t!�ǿyXAm�� ��<��]��i�"�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\蟖�S� ?�0��E|�,°������R�wX��r7�r��#[�$ԠI�*׿j�h�<�1#��Z�����XP���ct�:��RE�QS����>�[�W���ѥ��e�c�dט�w����j����r�C�M$�1#��Z�����XP���h�5,Wl�/�O'�=��Z������p�m~|���u�Y���\1�Z���=�Ln��S�W�7����KPy]/�qF��$�9	��NNT!�5_~\C�~��/(�����@�{���ĠЋ�l�T�Q��O�بeD�I�1#��Z�����XP���#���1���Q��ǺΕ�|7J���UĈO�����vޫ��%�%����=�ܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L':�N�y�w��ݪ��°������R�wX��r7�r��#[�f����0+W���F�^��NP�b9������U.6��̞��>�����Dɵ�p�AJ�e�$�,W��+�Ds�`��=i���Կ,��_Vl�A.;��L�O����K��5����`K�z~~�Y_" �g8Yw�H�MPq6.JHn��z������h_ъY�7#�xIQK*QYc����it	�T$x�����
iEE�G�����zP�����1#��Z�����XP������0/�e��9�S��8�U]k�(���B����_T���a�aq���U�n;p�m~|�֙X�D��U9����u�I���'����=���a�>�*�).zVW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�pl� �PP��ƿ�c �B�dH�7DR�i�Ρ��˧T������X�p0�&�����Q�a5���nXZjwi�U���Mչ�����Y��n�Z(Ρ����u�PBxN��X*d��Uf�Y9��_QzMy㥁�hK�'�njVfV)~�`V%'�\�*�c��i�#uA��I��'��b��v݋N�����[���S��IÙ=�H��"~6���aq��͹��e�[�.ᬵy����`x�AqeGfB�.W���ۗ'!�b9��!�`�(i3�E����FZ鎬������_�,���ܛk��md���{�!�`�(i3���+�J��Y�{'%s�6F���y�踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ]�N��&��v1a{J�4��pBy�p8�(�E?�o>������
��M����A�m�([}�@��L}�
�?��e�S��@��Vd�����<7u�r�&Ɓ>i[�ͧ�?Y�f�kN�ı*�7`����\Z��K��4����/�����N���Q��B%��>&ޝ����9OS���|��{�r1��j��M<�DO�)�U����I���
�CӞD���:�#�.��N�x%�4�.rM�1.ZVRѿUJC���d��ݷ���r�)p�ȷ��}�
�?��V5VM�d�bc�-d_�k�:A�	S�r��AR1<��J�@Ym��`�z��Y��),�B۸�1��6iRl�i3�ki�a����0��4�7��r��]�N��&��L�t��n|�%�|>��A3�(N��㎏qló]�b)�L�uf�Nd+l�Yҽ֗��i�ܰAb!��u�ϟ��7�4"���(h�:��
��D&e�2l��4(�de�QV踫g(�r�N�ǁ�f�TpD��ZOU����q�f@ ��*���v��W5���i�0�OgA�I�y�?ܔp�l
d�R�.��On��M���I�m�J�!�L�wV�}�
�?�a���k�_�~v� 1����/y��g�'b�t	�U���C��O]r�<Uee��~j�������I7��-5r�p =(�a(􆿳���2����.vے�(�i�p�� �&�K��5��]�!��M8���	D%��_�ͅ��I4��欱���j����թ�g�8Vct�:��RE��W��_�ړ8���/����,D�
�t�J8�=��ծ��:�a��Y�{'%s�[�&B�踫g(�r�N�ǁ�f�TIX����%V�����F˯�+)�"j���b7|#9���aZ��qA�E,Q�\C䗣��S_�����+�J��Y�{'%s��.|Z���I7��-5r�p =(�a(􆿳���2����.0��jOT���b�S]�I�$� X�]�!����w�Հ��A�YHm�QXv�5���f�g���Z�!K��tf��
_�n�@/%{�;����f�kN�ı��U��+�Xa�H(�˕-+��B�G����n9�}������ݼ��s�G�7s�9���on�-�6��
�jW��D���M���o�G�m�?%^�����I7��-5r�p =(�a(􆿳�ټ*w2�56ݓ��E�/�������� �mDƇBHx\�'���Xw s4S�'�i��`�z����k!�\Z��K��(Ko�yؿ;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J��H����� �����p՚��l��Hr�<Uee���R�}vJ^�k��76����,DTc�~y��i����u_7s�9���on�-�6��
�jW��D���M���o�G�m�?�{|*�"�Vx�%L��W��_�ړ8���/����,DTc�~y��i���n���g�p8�(�E{p7�j�pܔp�l
d�R�.��On��M���o�G�m�?H�OM��`�<'C�q��M#��W�s+��6�.6+�ii
��U�e�7����	N^�U{xN��i>r�<Uee��H�ʱˡj�:�IL���,D��=����;��krk���:�a��Y�{'%s�[�&B�踫g(�r�2������"�*o�yG�qڒH[91�Z���=��L;Л��|#9���aZ��qA�E�푧)����������H>+�w��0z�cUL�n����4����it	�TU����z~���ӯIJ ��`y���h}Nw���eZ���08:�}v����]�!��	Ǹ�y85��L�@��f����k��$a(􆿳���2����.\�#$�ÙA;��W���n`5�fK�\w��0]b!��u��չ���1�JS���$�q���U�h}Nw���\X��!���t�5�AԢ�a\��F�dHS�`�\��g()��ikp���H����HRCJ��<om��ڱ{a�ܸ�8���/����,D\X��!��Ot+�z��AԢ�a\��F�dH�i�rJ�(�g��U-�e,%�0g��Յ�HN9�5���u�L�xZ��j�
�iB{�Z�_�vW4��`��Q��ǺΕR��ӟ-�F`���G���`y����@����gGf���ѩj�T]t��T%ٝ�b�Bϱ���w�K�1c+����Y~�y����u{ᵿ�����"X��[��Q[R�7�׎o�|䖬n����U,�(�)8���0y�	��sC��#���FӪ�c�g<�g��U-�e,%�0g���Y�l��u$�5���u�L�xZ��j�
�iB{�Z�_�M�l��S�J*�Rs�08�b(������#oM���Øf}�
�?�����}�)r����'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,D�=P��[��1�U���]�!��	Ǹ�y85��L�@��f����k��$A�h��+Fen����9��0|~�LL�a(􆿳���2����.\�#$�ÙA�B�r���n`5�fK�\w��0]b!��u��4�	��������Oˊ��C���g��U-�e,%�0g���b02�O(�`ʂ�7s�9���o>��l%i�-�u��Y'GU�_V�"��Q]� _ό���.�}�
�?��G`B� зq8�Ј'���Xw���,DH�v�����] 1�0µ�]�!����w�Հ�*��9W��}�bo{W7s�9���o>��l%i�-ݓ��E���p��b����b�g�Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/�I����"�CeFJ5x�_�k]m��D+_{6��lJ��튝�b�Bϱ���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X�v1a{J�&��	�>�y��Fp����f���,(���B����: ��ao.\C�kHgN�����`y����@����gGQ��6��'��o\�B/M����*����^.�]�|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�j�W����+G��ܐƇ:Vxp�ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_S⏸[��!�`�(i3��lJ��튝�b�Bϱ��ᵉ3��鑘2����.�>��왩�/s�1��p!�`�(i3"�,�>E��P"G�wk�١��	;q���z
A��Φ�gz(AٸI))����A�m�(��A`���*�8���/����,D����y�[�l��姹� �Xz���úAV�!s���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�[��m�U����#3P��I�q��T�ٮ|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�����bp�WdM4@ȴd�?�V�^!�`�(i3xZ��j�
�&�j��1�a-���7a
��r��L;Л��|#9���b!��u�[��m�U�H"҆>X�����鰲�O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g���j�|�{'�v1a{J�j�f�At��usR+��f���,(���B����: ��ao.\C�kHgN�����`y����@����gG��l��`��Ĵ��ޯiڡ�F1�4W����㞮|�,
���]�x}NI0���ԏ�.fOe	��q��"o��I/J}�
�?�3�:���E@m>r
��1�#��d_�k�XLF�iB{�Z�_��׉p'*EF���L��b��v݋N�����B�d��,	.��`y����x�6�u�Xݫ,��G!�`�(i3!�`�(i3зq8�ЈF&|S���T�\ ���&�����~��U�*�şxˏ1�iA'R�	�yvc�]k��lJ��튝�b�Bϱ�����7���{r��'6���;8=�g��U-�ez�r�6�>��왩��k]m��������fQ��Υ�d[gȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g���j�|�{'�v1a{J���!<����㞣ɐa�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀ*�şxˏ1��o\�B/���2�>�E����FAԢ�a\�D�����R�`�|��K�z�!��(��-<�'++�g��U-�e,%�0g���j�|�{'�v1a{J���!<�;Ai�ŐP"G�wk��r)��ׁ�a\Y����)���8˩��F�{a(􆿳�ټ*w2�56d�x� �q5=��)Q��E����FAԢ�a\��F�dHw(��ES���v�8:�x�3�Aga(􆿳���2����.〧I���}�Z'BY��lJ��튝�b�Bϱ�a(􆿳���2����.〧I����뒒�����lJ��튝�b�Bϱ��f8�;ʄ6���n6�R�wX��}�
�?����D)��C�V���3�ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀ�6�S2vTDZ��O$ғ�vq���q�41&q^�`
�c��><�$��;mQ��8���/�I����"�CeFJ5x�_�k]m����DބiMғ�vq�\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gGQ��6��'Rm�㭼�S}�S����=�?I®|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�G9�:Q����Z$�x�߃`úC�P"G�wk�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.JL���Z'#y�>�)L�����/s=s�^�?�/S	��1���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀCeFJ5x�_�k]m����\�6��dR�8/\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gGQ��6��'A�{�>�� ��
tCtHC�'Ϯ|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�}c��ko#�/��y?�-� n���a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀ�6�S2v}�k�����|	�WIғ�vq���q�41&q^�`
�c��><�$�X~��\��o����׋��`y����@����gG,#�g��C�x!�H�M>��#GK'q��T�ٮ|�,
���]�x}NI0���ԏ�.fOe	m���h��D�P�E6���2����.0��jOT��.m��K�+���w�Ѥ����f���,(���B����: ��ao.\C�k�ף�D�~R��v	�R�wX��}�
�?�G��-�HG(�b�'Be΁�a�n��xZ��j�
�&�j��1�a-���7a
��r����~v����"X��[�d�a�4$�b!��u��Ɔ ���Ve��˅�q��T�ٛGS�����n���㬺ƃ
ᾆ�x�T�\ ��i3�|)sՀ�Oi9L�:�k]m����lJ��튝�b�Bϱ��R<�����á�~O��L;Л�����Øf}�
�?��I�_Pg<�%��g:�����<�ׅ��A5W��v�8:���h�|!\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?��I�_Pg<�l��姹�n4'����3
�v�v-}�	mp���g�<)\[$Q��
�̞��>��b��v݋N��������(($��R�wX�ո@����gG����<��y�@�vFn�H�~M�!�`�(i3!�`�(i3!�`�(i3!�`�(i3O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv���9$��i�Yi䚠疛!wFii��.�m���!�`�(i3!�`�(i3úAV�!s���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u���a�vw����~m�(��k8w��?L�@���wp>�\�H��/SggR��N�$��a�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X&U;��]�x�'��x!5����z�Ji�!�`�(i3!�`�(i3!�`�(i3�k�XLF�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'؁C�*&#�4?�o�5�h�B� ި�6v ӫ/��m�h��"��зq8�Ј\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?�rS����u�}�Q���GM�о٫�S��wE\�!�`�(i3!�`�(i3!�`�(i3ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_c(H޵D7W�:����p�A�z;#o"�I0���ԏc�r�(������^.�]�|�,
���]�x}NI0���ԏ�.fOe	��q��"o�d�a�4$�b!��u��V3����C��z���2=��h��f���,(���B����: ��ao.\C�kHgN�����`y����@����gGQ��6��'�֤���n���6����?��ө%�Sg()��ikp���H���ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����]�gv���J����0;�����5u�q��	�����aq��3���WQ��|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�G9�:Q��F��P�?��4�+��_��A5W��v�8:�;��so��f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/����,D��ǉã1X�v1a{J�Bz��s�V�c���,NY|VO�⅘��a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀ�1r����Ɔ ���Ve��˅���ө%�Sg()��ikp���H���O�=�ͦ�١��	;qS�>�!/�_�n�To�[r��}k:�>�hy��T�\ ������q�f@�]�gv����U�h�ݭ$;�
��f|m�(��k8�k�XLF�iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��!&��F�!�`�(i3!�`�(i3���aR�}�
�?��I�_Pg<˃�B�1Yw�Yi䚠疛!wFii�?�(�L��>�f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/�M��%�p@!�`�(i3J�W��7/�CeFJ5x�_)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��cP��N�3��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����]�gv��L_v,<=��}�I���Fn�H�~M�úAV�!s���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�Г�����!�`�(i3!�`�(i3J�W��7/�CeFJ5x�_��\�6��#P��Ѐ�5�h�B��ME�R�, �EM�3� �a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ���sC���XaZ��qA�E��ǉã1XBz��s�V�r�G� Y� {l��	[�������a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ���sC���X!�`�(i3�@����gG���y����7B��[�<?Ә�%"Q�ܦfM� �in5�҇�?����XzR+0��^O�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���%^���\����iW5���(�xW�A�&hH\l0��F��j�mV��5f�l�I�SCp~z�r,o �#^{���y����b�Ա,G���P��w�T:~m�iX���]�aq��(ք��h��Օ��qvdЧ^{�jt��zh+�,�l��=5;.�����/�q
�@�#��fx'v�ao.\C�k[�(��PJTXO�[?v���N���.('�?��&^���:�����
��PР?�:7.N�ӃHoh�:����K M2f�����������ĬM$2�à�Z��ޛ_�.�˨/MKo����\�R���	��}�
�?�Q١Ӿ�$/s�1��p�E����FAԢ�a\��F�dH��e@�N�] �v"��x�l�<Ң�8���/����,D'���+)'J���|�b1�#��d_xZ��j�
�iB{�Z�_��?� Zh�R?�R��nI4�p� ^�b��v݋N�����~DJ��/�a(􆿳���2����.�E ����$,K�9+�/���p�������������B��èVϟ��7�4�I�N$Z)ݝOv%F�YCs��$2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�*���
Cz�%�+Z�\�1�O��k��`Zo�(:�J��(q�8�(��y��ڲ�ؠ�:�f�Nd+l�Yҽ֗�G��e��;��|B����Uk�������	}�@���F����N�ǁ�f�TIX������bT2�5�O�%E#PY�4Eb��Y{�o��e:-�t�sH�g��6�e4����b��T�Q5�:�2� _|�8U�.@����J���?'drD.A�s���Z�y��J�\�=6�C�&���	M��3
�v�v-}�	mpB(p`D҉�Y~�y����u{ᵿ����?ڄ��5�O�%E#P.�`��ai�}#�U��*��Y��!�`�(i3!�`�(i3W���y�N�#�r��8�GQ����'V�Ո��+5�4��c �&A�5I��RhF�� ��*�C� #�~	�D�t�3����%�toqP�N�ǁ�f�T�A(夽��׉�/fI��)���W�w��fDK��l���V��J��n�f_���� � �k�3|���x��@��ǀ�D=�A���ۖ��S�<Ԣ�G�nJ `G�p�P��n7�_@;��|B���r�����Ͱ�Ǭ�j([�NI�P�6���ퟓ���2�b{��3x�В&=�y�q}��#VL�^^J��n	l��Q;�im��ȍry��	�D:���@���k��!�`�(i3�F�7��Y�
�cc�V��ݚ�Н�$Q
ˋ!E\1�1�ҕ-��3�^�P�qjhbvk~�#x6�V���	�Y~�y����u{ᵿ���$o#[�L\!�`�(i3^P��:w0I� X�1���Õv��9e��/�7�!�`�(i3�2*Q=F�k�mD#V��A��`-!�`�(i3�po守�ud;��,4��V�;e���`���ҕH{6��!�W��!�`�(i3�
ۼ����F#I�%�[<c�=,!�`�(i3�O�G?X2�K��2WI'�=��y�ݚ�Н���+qѭ�+g[�!�`�(i3�M�g����H��bf�?ǉ�=�y��j��k
e�3+{�i�m�T��!�`�(i3�6[��u�9k�\,���m�
��,!!�`�(i3扈�s.�֡mh�l�Rk�X�
�s�!�`�(i3p�n���:��]]t�GR�D^�6hg�}��wӨj]h���6�ü��k>B2�2�,�^Ȼb�8�dX��3x�В&=�y�q}��#VL�^^J��n	l��Q;�im��ȍry��	�D:���@���k��!�`�(i3�F�7��Y�
�cc�V��ݚ�Н�$Q
ˋ!E\1�1�ҕ-��3�^�P�qjhbvk~�#x6�V���	�Y~�y����u{ᵿ���$o#[�L\!�`�(i3^P��:w0I� X�1���Õv��9e��/�7�!�`�(i3�2*Q=F�k�mD#V��A��`-!�`�(i3�po守�ud;��,4��V�;e���`���ҕH{6��!�W��!�`�(i3�
ۼ����F#I�%�[<c�=,!�`�(i3�O�G?X2�K��2WI'�=��y�ݚ�Н���+qѭ�+g[�!�`�(i3�M�g����H��bf�?ǉ�=�y��j��k
e�3+{�i�m�T��!�`�(i3�6[��u�9k�\,���m�
��,!!�`�(i3扈�s.�֡mh�l�Rk�X�Q��ǺΕ�A�m�(慧��a�f�?ǉ�=�2��}���zgm##��V5VM�d�4�|W-���Y��),�B۸��1(%"{����%>�rG6j�"Hs,/A�|[^�Vj�Ra�mR����
w̅�_��̶I�?g�f��Qө}�_g�?�H���w�1��YO�.Ŏ����%kR��������֢&@��&Zt%��m&<9U:����VK�5��&q^�`
�c��><�$���E��!�`�(i3ct�:��REvє�&���ct�:��RE3z%�u�܆!�`�(i3Ĉ���rl�خd���!sH�\!�`�(i3C��[�����p��@LC��[���Ը��q���đ_�������� "5�]!�`�(i3Y��'�����0��"��S8�TkF����v1a{J�Ώ�y�JT�f�?ǉ�=|�\m��sG���MY�{'%s���F����:�#�|$.@L�`�ui�Tc�!�`�(i3��
���;�r�=k�Hg��iqk�f�?ǉ�=q�\E��0���N��t�3�����D� ���!�`�(i3u�l�T.��:��]]t�L�t��n��Q� ��!�`�(i34]:C�2Y(���˜V�
�sǟB�'��a���r�N��(�����/��@��e:$h�7�cl.�	�C�!�`�(i3�Q}mҁ�t����sM�yx�,�G�1�ix�b�8�dX�↨q�©�����<��p����Գ�9�^N-����Lt�iZ]XF�hx��G��!�`�(i3 k��v(�Âv����Y���a\Y����+���LQ�f�?ǉ�=�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=j:�Mpp�}�(�-lc4�j
Թf�?ǉ�=��X�u��
)\Y����4MT2g�ȨQ�?�Q!�`�(i3���ȍry��	SƏw0��П�+�
8'���Xw�j�7��9*�"FP>���뭟Q��ǺΕ�A�m�(�]�	��B7Ԅ��SƏw0�����.>H'���Xw�j�7��9*�"FP�jV�$d,H�Q��ǺΕ�A�m�(�]�	��+#Cxz!B��2��}��̏A��?�ϟ��7�4Ï�6]S*�N�ǁ�f�TpD��ZOU	XT�1�wӨj]h�z��?�9��V5VM�dn�0�I4��欱���j����,X�|H*!�`�(i3u�l�T.��:��]]t�L�t��n=蛗�+N���������$��+#Cxz!B�`
 ֢����oC���b�J
�g��*�7`����\Z��K���䈷UJ!�`�(i30q���Q�L��!�`�(i3bs��2[������	�;�ݚ�Н��\�LtF�/�X�h��E�i�m}66j�"Hs��ˑ1Ms�����x����A@�Q��ǺΕ�A�m�(jj�*y��}�+�ϸ�i$x���z*�7`����\Z��K������]NS��.�g3Z�j5�{�ݢ��e��[њl����{O��c_`J��Y��)�.����ߤ��/��5�O�%E#PP���x�NS`|.^~�/W�/�#+*f�GR�D^�-�����6j�"Hs��埏���7�VL%�ǅ�����xF�~B�@o��[ea�8��������?9|[�,HJ
 )�1��kV��o5]�Q;�im��ȍry��	3A��g�5���9dss2����`�|��K�z�!��(��?�&xHC�Wn����������\����>'���������6%�a�]{��_G�D�� ��ۋ�/�ͪ`�3J�V����U����\��,&߰��U���BA�IH���O,8����������2���]�!��	Ǹ�y85��U�z����@{2귑��?4��44�~[ی3�ASƏw0�����.>H'���Xw�j�7��9*�"FP��� �mD�^��x�dŠ�Ŋq�\E��0�aR�J�}#�U�����Y)N������	\k�`��B7Ԅ��3�kM�}��s.�֡m�\�&e���Q��ǺΕ�A�m�(It8Z�QCf�?ǉ�=�!�'
k;r�=k�Hg��	��+@f�Nd+l�Yҽ֗��J~xAU�"VA�ڦ�c4��3vS�vN��%u��f�Nd+l�Yҽ֗��J~xAU�"��=����t��r�N��(�������0�&�ͭt�%�Z?��<�ry^��Q}mҁ�t����sT��{B�z��z6Y��9$��i�B�@o��[ea�8��������?9|[�,HJ
 )�1��kV��o5]�Q;�im��ȍry��	3A��g�5���9dss2����`�|��K�z�!��(��?�&xHC�Wn����������\����>'���������6%�a�]{��_G�D�� ��ۋ�/�ͪ`�3J�V����U����\��,&߰��U���BA�IH���O,8����������2���]�!��	Ǹ�y85��U�z����@{2귑��?4��44��+�5VlSƏw0�����.>H'���Xw�j�7��9*�"FP��� �mD�^���ިMiT�zq�\E��0�aR�J�}#�U�����Y)N�����:�bC�t�{#	�x�z��?�9��V5VM�dn�0�I4��欱���j���֬���[pq�\E��0�D�0���t�3����%�toqP�N�ǁ�f�TIX����+#Cxz!B��Aɀ��	{⟰�&�U���H^�N�����:�bC���=����t��r�N��(�������0�&�ͭt�%�Z?��<�ry^��Q}mҁ�t����s2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha�Ko��m�\��5/<�KǣDޛ_�.��)n�w�'��Lk}t��]`�L�FZ�1ǿ��^Ý���z4x��x�L�FZ�1�M�ŗ\�'	�?��[Q��Ш�^v��[6"�I�?g�f �H�Z��1]���%ӳ3z�]��t�iZ]XF�hx��G��!�`�(i3n!��i+�ť�n8���L��g�I��RhF��8usl�z ��ݚ�Н�w¹��<d�Ji�];���w¹��<d�,��L���?�Ho2��O%��<��=�>�t����oD�c=p�J��w x�·���~X�~���$^!�X;p`�����?�dv��oTN֢&@��&��|��p8=�[Ǵ��p���@Z�_F�k-�H��bf�?ǉ�=�|�)՜�4z�Gb��P�!�`�(i3|w�{P^K���3�<�p�� �&���ç�A!�`�(i3�\�!wn�ř�3�<�p�� �&�J�I�'!�`�(i3+�uB;y�3�<F��׿]!�N��y|N�F?P�.!w�E�U�P�)>�
��`�;��%YM�	�v�3�N�ǁ�f�TIX�����^�̷ؠJ��:����_$U���b.����{�vWދ�qc:`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��a���k�_g��������B���+�ϸ�i]T�o8�'��$zө���)󷥯��v
*J�X�$���jh��f�+�t�3���D��m���*�7`����\Z��K���&����$�HN��R��?�d���&��_$U���0�(j��0o�{E}́�9��,'6�F��K�J���1&NXs���ls�uH��q�/���˚����Z��L�{	����F��׿]�v����D�ه4�tZz_nÑ2hꬺ��1�$r�t�}iV��	��y�� �P�qN,t8��og���;_��8W�w��fDbYގEV�9^�o�a�!�`�(i3��;_��8W�w��fD�M߯�Px��|�������x���	R�N~)�j��N�����?�d���&��8�E�"0���a?�5��	}�@�r�<Uee�N�����$��̼�K���Z��L�{	����F��׿]�  ����'Z鎬�������(���[���-��G���۵z �+5�4��c5 H��d��$Ι��o���ls�u!27Ք.+��o������	fd�c�=���L�:w��G$��a��V�K=�u��HN��R��?�d���&��@��i�fKw�R���y��0�J���y�(�\tu2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڧQ����7��� -Q�7�p�D]Ї'G�+R���o��_�Rv�䩲$��8��I�:Fa�7���z��O��Y#&����"sS<�0�zG�������&G;�x'_|~�뽢�7;��1��J�b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-����Dw\����>�lj�Ǎ0Y�{'%s��v�9˞�g��+˘\59:��lJ���l�}0���	��+@f�Nd+l�Yҽ֗��
i#�"��$Ι��o���ls�uGR�	A�"HN��R��bP�63Z�t�5ߧE4��Fr��j������"��Q�JL����	ǜ�N>$m<m��ʘ['Ӭ��yb5]��o�������Z��@?d�s�8K,Q�\C�8�Hj\���n��\��d�٣��c�A�L'�c�Z;�b�R�wX��d=��¾ȼ���4ܱ�������{(z�Sb�f՛ةmy�m���~��Z���Rk��4�����b	��}���Z���7߷M�,���9�ԖY]�蒾�$O�L~�4��>m~�jxBQ%d"Y�9��$9��ճB*�2����CbZ�� Le=mlf�u�c�n��X�L�5_$�՗�(�[�#}�P)-]��h4W�7���\��	���.��yV�$�DK{Eȷ	{�z�� `�*�bn���==g�׷kM�#�> _;��i�1�CɀU��ڞ���ˇ���/�����P��?�N�ޖзu��v�<fGeY�:[d�d���̖b�K/P=<>|�`��c5�J��0�~�G��-�HG($R�i�Yl-����<&Ѳh��N�M��n��mC���!��1{�F}���V6��}�.�p�'�B��?+���נ2�9��V�9!�`�(i3!�`�(i3!�`�(i3̓@?5����T���b�Bϱ�� Q`)��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3/��kOT�)�����m�q�/�Wv�A���U��)���Y;e�iK!���d.O.C�U��B��-����A�;�>��z����8�Hj\�����1:��xjzӝ���I(͂��-����Dw\�����b�S]���o"83�� P�jc�8�Hj\���M7#� �6���n6��dh_��tCdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3G��-�HG($R�i�Yl-ۼ��%�ۙ�b�S]���o"83�C�
���W����Uh1݇S��;�q�Y{�<���^�[�-l��NMm�P˙��b��Bg�Pڹ�ԑ�b�������`y����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끓��~�L ��j�Y{�<����
�9�v�T�T�y�8�Hj\����Fl��m�q�/���e���W�ɸ}(��:)�
�9LeQp�K���&�K�VF�P����9��g�ܧ*ys@B�u�.��.f���s��1�y�n�F�:)�
�9o¶D�ν��jd�	�!�`�(i3!�`�(i3!�`�(i3��j�4�q��_N��¼��=B��u��;���� ���J���*j�B3L���(�Q8;��|B���r�����EHd
0Ki�|2;$�J��7�OT�,��7=���bڕI��.Eqb	��G��W+��W��P����9��g�ܧ*y&tS�D������_�t���׻�fĉ>99��;��|B���J������
H=V��	��y��%����,$�R��aT��3G?�d���&��ҕn�s�[dv�*s?���[`Cw�H���-k��O�)"���.>mT�Ɍ-';��|B�S��sF����b�S]q�6��^�!�`�(i3!�`�(i3��$�\%eK��J�x"V}�IUr��� �&A�5e�J�Pn\�pD��ZOU�S��;�q뽢�7;6ik!�S���{ �4"-�"#+p:wH��|2;$�JأͽgF"?��7=���bڕI��.Eqb	��G��W+��W��>�:| ��k�4eYy�tDWfD.v��W5�!�w(�y?w�R���y�-.�zP&K��Q�m��)� �.�g3Z��~H?��2�.�|�e$S�Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h^·ʌ�C��]���Ҙ�9 �/����P�����
T+Fb%��C��:O�����=�w�����5�O�%E#Py�y�Ż�"�_�0��(����5�?�J�Ń��ɖ�2i�螘c&#VL�^^J����S���� "5�]ޥ0D��/��=��K���0P��h�5,Wl�/�O'�=��hQ�GvESƏw0�������_�H�f�M�&�;^�6#9��u��n��ݚ�Н����Y�l, 	�I��0��:|z:;�<%�a���(��	YRF!�`�(i3ct�:��REa��ZAδ��כ��p�,��L����+�t2�0�趦���o�Hc�U0�!sH�\`�3J�V����U���@��������=��܄�H#�"8��!�`�(i3;���[���{s�ܱ?'�=|-�e1|E�A�2�1#V���<�dv��oTN֢&@��&���Mڷ�21!t*x�S.!ū�ez��k]m��,�۞��	�rVu,� �{k�h�+|�c�$�t�]�;���VС���u_�P�v	��YY��
�iC>N0Θ��ݚ�Н�bs��2[������	�;�ݚ�Н��Q}mҁ�t����sX� �Ĭ1���$L�9���3v��u� 
~�F�,���XF:����k!�\Z��K���^�̷ؠJ��:����|��Li���Ay[����=ME8q��ǵc�;-;*�7���d5z�R��T�\ ��;��|B���r�����Ɔ �����Vd�*J�X�$���RW����C�x!�H�J=�m �T#��(�&�.�g3ZrZ�0m�\�9�Z�y�6��s
!��QS��:Z�����n!�'��iF=�xo�R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G�dE�h���|f��ӡ`��R������s��ꬺ��1�$r�t�}iV��	��y�� �P�qN+M�ᴰ`��~���.�;��|B���0�2u��$L�9䮏��5���%��;_��8W�w��fD���}l�g`���U��t�i��˦���X��lM�Ҡ�N�����?�d���&�C#/<���q�*���Nj�MC�%`zI\��!��6j�"Hs����]��.��M!��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�i"����X��d��9�>�:| �II���؄m��+��jTʱ�8F0_H��w�Sjs���V��o5]�Q;�im��ȍry��	��M����3��~ �X;p`�f�Nd+lJ�VeSZ3&�=�<α2
��j1dM4�<"NU�:|��6/��������рӚx�f�?ǉ�=R�c4!`���������+��c_�B&��p��Z�%P{�W���`moF˯�+)ƍ�����)ύ^��Ĉ��r�]@�����ՔiyV�[R�^Ƒ��!�`�(i3��4��#o��
�cc�V�����b�y]/�qF�B�wj$g��ߐ�*׿j�h�<��k�+9=NM(�n��1�Z���=��m�B��dVkLs��dJ�+���LQ�f�?ǉ�=gR� �ұ!�`�(i3�Y�M���˻��0y��<0��s���4@Q�/��y��j��k�lԇ�-{�t�%�Z?��<�ry^�h�'f R�苇��Fe#OOJd֯�|�)՜�4�X;p`�YmC,iguEOJ�uxm�3���w�@V�?ZFw�N}�IUr��ӭ�
:&��5��=����t 7�J�[�_�C�6%�W��|K:�2�O
�� t�{#	�x�jsrCm�kz�6�j=j�3Y����/�sL���S��-X� �Ĭ1�e����:�ԑ�*V�D2U4��\w��˪?�-C
2��>�q;Rm�5�O�%E#P1h#��x�3>�G5��,vQQA�q�m�,~s����2���ܝMM
��,=?�d���&�t�{#	�x�}������ݼ��s�G���>�9��l�?3X�`���%]]��ToHA �I��)���W�w��fDv���k�#?
]w<�9w55^Ftw⪞mf��j�Txk^�a���~6�z�����ϲ��Vo[���˚����Z��m�����G�N�*J�X�$�@�J��L�jA��|�qG�U�I��O0Y�6j�"Hs�ĖYS⪞mf��aT��3G?�d���&�zY]�埅4`v�;w6%���7�J-I�p��g���y[J3�j\{ف(�7���<��Y����}J�|���|���>�q;Rm�5�O�%E#P1h#����5��������o��D[�h��4o�ݪ��H��q�/���˚����Z�׽F,���s+��6�.�Rhy�$�������;��krk��ꬺ��1�$r�t�}iV��	��y�� �P�qNp����*aT��3G?�d���&�zY]�埅�t�į���W�\m32�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��iڈ(���iW����u7B�k"-�� ���J2��������������]9�(b���J��:����Cvu#��I�?g�f �H�Z����dn��A\^�N���������%kR��������֢&@��&��k���t����~�.O9��Q��Q��O�بeD�I��k�+9=�]V�H7'�R�^Ƒ��X&|a�#���8��'W�Ty��5!�`�(i3���0/�e��9�Sw�%b��G����p�><��d5�:�w�+���LQ�f�?ǉ�=�ܼ�Y�{ �=�%�vє�&������0/ܤ�(g��V(�G�&���k��,�:�N�*�x֭�h��Oo��0��7�˺�Q���f�?ǉ�=�M�g�����X;p`�(���������!�`�(i3z�Gb��P�!�`�(i3�<��>��%@��4���~��rͤ;��krk��C\�2x���?V��j�c�[N�&ѐ�1Ʌ�Mi�������F�����7bYގEV�tպ� ��q_҂T�q�w���Q��O�بeD�Iѐ�Xr��,��d���!i�&+�eo$��Y�C|P���=MED[�h��4o�ݪ��H��q�/���˚����Z��k��u����f
t斃����u_z���]�D�ߌ�LM�a$���|f���s	��e�.�g3ZrZ�0m�\���ٕ��ж���X�*V��	��yG��Γf��Bp����̳Ƒ��EQw�R���y"O���%jm
����+
o>�I�	���j�[;���M���R'),��`�ka�9ϥ��;��|B/B�Â����dn��A�9�2�L��f
t斃|�q�^"��.�g3ZB�ek�5W�Y��N2H���/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ����s���BK9r��B+��d�<��I�?g�f�,�� zr����$l2�W�K��V��o5]�Q;�im��ȍry��	w¹��<d���<
DN��$wq����+W���F�^�Y�7#�xI���E�����o)�]rH����8���f��9
���M���R��ӟ-����6%�a��Nm�ju�|`��P��a݃�j��C�`�/�t���E���� ������O�z���5$�<w����0)]��w�b^X�P��EގV�ڇ��t��˳3[�u8����ꀍ�@;w�$C,0�?����_F�k-�!�`�(i3���*[UxG���%>�rG�B�r�݇a�/!O�$-q�0c$�Zt%��m&<���_L�b�����Ee[u�;0�f�?ǉ�=r�x�e�X�k��rݾ(����C���h���?V��j�c�[N�&ѐǂ��%D�$o��)�ͳ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���L���Ŗ6$\K��p�>&�+���LQ�����_��j��N�֞q˩���.|�YtA[���Ŗ6$\K��&b���E�vL������ur]p�+#���&�x�.E�FY��+c��8���ݔf�zE�񪣘yg�U�։�������� h9�=�^�a�	�ӪЪ�S>f}f�Y\%wj�j2�%�}W���8�=�w�����5�O�%E#P��_Ѭ�Q�vC��Mi�ʷ��A�21�ri��WH�1�:�Ω��maC�S�s8���\���PM�^-q�x�l��1:�N�*�x��
[N<p�U��֜��3�X;p`�Q�%�+2�j;��q,�?�Ho2��ݪ��t����$�fC` ��\�H�MPq6.����gQ'�|ݔ�3�(n�'�f�?ǉ�=$(��>��������	���i$;��|��T�.�l�.θ��q����k��,�:�N�*�x3Lv	̅���X;p`�(�����֭�h��O5�tx\s�l.�	�C�
�:qEp��:��Z)�"r��^&���贵[�л���7#���=
 �4���ߩ��ݚ�Н�p�n���d�)bU��� �Y.�.�g3Z�7�4��~��=�>�:|]η��E�<���5[�������0j|�~{b62�tstJ��:����s͟;)f���d�jO)īIX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�+��%�k<a�E�Rq���my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н��}�АR�38v�s3~�0�����&G!�`�(i3+��%�k<����m��5vȹ|b�7�ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��@qz�_vrrL�����^�%�P�m�V��	��y�f�HYs��uF��82�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0����t��[���P��EC�`�/�t�KV*�3?�|��T�5�d�,W�He�!� U����z~/�}��j,NJ��:����8���SY�N�o��C�0�_E,�8�o��_�Rv�䩲$��GQЌJ
�յ[+8����"sS<�0�zG�������&G�wӨj]h�(%����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩ�-��)'�E��ȷ��#o�]�ʄǾH/�d��_�mS8<�n�ݚ�Н���4�*BqC��~�;ϔW򻐗�NGq���ÌZ>u�,R�� h�ҩ��wӨj]h�(%����+�uB;y���O�	���lC��U�T�\ ���:5A��pfĉ>99��A0ok�ª���l��������t�|ݔ�3�5�}�]�����nv��~���$r@H�RtV�^;�jmT�#��|�!�[�w/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=��,�����!���2�(+�uB;y���O�	������v�h��4y��ij��X� 2!�`�(i3>_�Bnˌw/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=�1�(�yj�!���2�(+�uB;y���O�	������v�h���ў�L��-����!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3�	��x��ݚ�Н�����l��q�P�oV4ʐ�}	�[���&�ŁHL�U���W�����&G!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1�B/���q%U����z~(����(]�U����z~)���	6�!�`�(i3�Ra])n#���r����!�`�(i3�� ߌ��̷_��yC��S8�>c��6/{v=~P0:Q+�3yK������v�h!M�T�ĥ��P�7� �:5A��p!�`�(i3���F��O��ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=�[�P�X;�Z��;_��8W�w��fD[�P�X;�Z<0)��TG䟳��LQ�%�+2��k��kK�I�Q4p�/Cj���C�1A%^�Q��U����z~/�}��j,NJ��:����8���SY�N�d�}����U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�{k�h�+E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l���{$����^V���!ֿ*Y��b"���LQ�/81tSjv��wӨj]h�(%����Z鎬�������(���[���-���W�6?��jsrCm�k#��2�bD�=�^݊��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M����m#p��ܸ2߆X�.�g3Z��S~����l�I�k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϓ'�al��p;��|BB�Q�ˇWv�A��=a��0� �Jeh|�*�7`����\Z��K��7�,�B/�Q{z�
wb����T�}ɻ*�7`����\Z��K�����6�~�5�O�%E#Pe�6&	 �|��k�|��SSB������a�v'�m����o��_�Rv�䩲$��GQЌJ
��`���φ��<�6�15���Dl=*�QN������"sS<�0�zG�������&G�0�9&،�j�W����+G��ܒ���7�_
�uz!:�X	��sC宸I))����A�m�(mq?��qU�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!C�� R�Q�&�2���)x�?{���x.�Knq��5+*��d�@���G�X���.��ġ��,��5+*��4br���qP�V>t'�̗�����F��~1tSjv��0�9&،�j�W����+G����v�9'�͘6��q���j�W����+G���|��nZ����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끣�os�鮊(=�"v��Iw�6!e�C�7ª6��J�����_�U*��ө%�Sg()��ikp���H����c���鿉�X+�kQ��v1a{J�i�\��ou#�m ޶&�hbvk~�#x��#�H�޼QE1��v1a{J�&���e�� տ�:
hbvk~�#xo�������Qטg�u2]c
j���l��姹��*�ɿ�4J*�Rs�08�b(���,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��LG9�:Q��Ĵ��ޯi�-Qq��Pn9a�Fc��Ǔ��K��v1a{J��blv�Bo��"~6���aq������n}L�I))����A�m�(�l���q�b��v݋N�������H��YTN��r8!�k]m��
ae���K���c����P7E����k]m��GTH�<�g()��ikp���H����7�����\�H��/Sg�w��'o����̜�I0���ԏ�.fOe	j�)6)-
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q��Ĵ��ޯi�-Qq��Pn�����G�v1a{J���!<�*Ha���J*�Rs�0��O�@�n�M?��h�k]m���E��Y��m���+)x�?{����}9��|�G9�:Q��Ĵ��ޯiڼ�ze��>տ�:
hbvk~�#x�<\��-��4�1���~!�`�(i3!�`�(i3!�`�(i3N��r8!�k]m���E��Y��m���+)x�?{��
0#`�1�������f�l��=5;�B�uʡ ޼QE1��v1a{J����%]+a�����G�v1a{J�&���e�� տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<�l��姹�n4'����3
�v�v-}�	mpJOv�����o\�B/u�:o+���	�����aq��c�:X��Wwl53�e�'{w#/ B!�`�(i3!�`�(i3!�`�(i3G9�:Q����v�z`���ө%�Sg()��ikp���H���R����� ӫ/��mt����� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�wbk�$�޹���M�,!hޖ�A$�P������5d�������y�:Fa�7���W"�P�K�0_f��3%�:��IY]��r$ɓǃl[�Ƶ�1tSjv� #��zG���J����(�u���p��,\���͔5��:m�\�H��/Sg�w��'o��Lͷw���]�x}NI0���ԏ�.fOe	�ߣ
����Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�g�s���������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��;�uO��Bu����aGl��Z����pG�p�P�$�c76u��r��M�yx�,�G#y�>�)L�Y�S�:3�g(���27:։�X+�kQ��v1a{J�c�Q$ a�3��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��uR�Y�A��-�R�͢��n-(�p��Kث��@�uj���V��H?Ә�%"Q䛚�z�Ji�!�`�(i3!�`�(i3!�`�(i3�I����~u͘6��q���j�W���]�B� �Q�ސ�՝.�&J�m�(��k8���0[�d�G`5[��{#Ÿ�&Sq�a"��ř�!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Ĵ��ޯi�^�0��ͅ�a��;���=����qFq�w�鎷�Z,����d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[�pI�
K�x�������E��0�Z�7W�:��G�z㤧{�̌�͚�3�_�n�To�[���9�P�4�D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�2���$H�WdM4@��z(�ﳔ$@PJ+5*�轓�A1�J�����)����Ҿm�(��k8���̜�I0���ԏ�.fOe	���X�a1p��j����Q�9�|`��Y�m�k?j!�`�(i3!�`�(i3!�`�(i3�a�x�]c
j���%��g:������	����^,�:��O�?�I))����A�m�(!|�α+���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~K�\7}�W, D�cg�}ŷ(K���}�;]MBg2Zr�G� Y�ҹnЭ:��#�@����ۭXX���E��O�;]MBg2Zr�G� Y!s!��xlJeYSWe^E˔ �y=kt��w��X����xQ�1���~!�`�(i3m��i�*�JeYSWe^E˔ �y=kAu5��ݞ<\�H��/Sg�w��'oD+���4Yʁ���Mյ��#�@����ۭXX���E��O�;]MBg2Zr�G� Y!s!��xlJeYSWe^E˔ �y=kt��w��X<���H1���~!�`�(i3m��i�*��9$��i�Yi䚠疛!wFii�v1[���b��v݋N�������(X��#�@����ۭXX�WŚl��E�d�G`5[��{#Ÿ�&Sq�a�"Ĝ���$��a�vw����~m�(��k8w��?L�@^?���W��j�[O����k$ !�`�(i3��䨘J�\mo5i,�Ĕi��)��ۺ��fyd�F�O����!�`�(i3!�`�(i3(*�O�q�@��i)&
�k�����oT`kz��9$��i�Yi䚠疛!wFii�1�В���,؁C�*&#�4?�o�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[B���v��؁C�*&#�4?�o�5�h�B�$5z&�D�� ި�6v ӫ/��m����	�����tj/�Ս��6Bj�!�`�(i3M�yx�,�G؁C�*&#�4?�o�5�h�B�$5z&�D�� ި�6v ӫ/��m���l]�f��EJ,�G7```+�ֶ������x�������E��0�Z�7W�:��G�z㤧{�r�(��mo5i,�Ĕi��)��ۺ��fyd�8]|Fl���1F#�֞q�F����&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N�����-
#?�QAmo5i,�Ĕi��)��ۺ��fyd�e�՝*U�޸I))����A�m�(^?����8������k$ !�`�(i3�~�7p����nt=:�+�_0c ���a�vw����~m�(��k8!�`�(i3!�`�(i3!�`�(i3׾ŞWsuz��"]c�#y�>�)L��H"҆>X�(JdT�ݙڈ�KK?B�&�_j�	�Ȗ@@��x�������E��0�Z�7W�:���p*�h<��I0���ԏc�r�(����I����~u��a�vw����~m�(��k8un��7� ӫ/��mt�����N��r8!c(H޵D7W�:����p�A�B��+ H!�`�(i3!�`�(i39a�Fc���M똡����o\�B/�u���a�x����r͖�k���$,�C�7ª6�JeYSWe^E˔ �y=k�2�u���e�՝*U�޸I))����A�m�(9�*��� c(H޵D7W�:����p�Ǎ�͚�3�_�n�To�[���9�P�4�D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�2���$H�WdM4@��_�U*Cw�Hm���9��N	{8G9�:Q��Ĵ��ޯi�3>٫F�?��"��II��jÇ+�_�n�To�[
MQ9�F�GM��QО��i/R�c� }!�`Uc�gC�!�`�(i3!�`�(i3!�`�(i3�a�x�]c
j���l��姹� �p�B���#;%%�.�4����
��\�H��/Sg�w��'o�֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@��_�U*Cw�Hm����a�vw����~m�(��k8�����9�Xy+�Mk��L

�F����&U;��]�x�'��x!5�kz���[h�b��v݋N�����-
#?�QAmo5i,�Ĕi��)���!D�����ӸI))����A�m�(^?���W��j�[O����k$ !�`�(i3��䨘J�\mo5i,�Ĕi��)���!D�����ӸI))����A�m�(!�`�(i3�����wP?��i/R�ce����� .����mo5i,�Ĕi��)���!D�����ӸI))����A�m�(�[?;$�\��E��0�Z�7W�:���p*�h<��I0���ԏ�?��Ds�-�w���+kGA��ݼ��r����!�`�(i3�o�5��!<��y�@�v�&Sq�a��z#׊;w�����f�l��=5;F5E�]q�hf��EJ,�G7```+�ֶ�����rS����u�}�Q���GM�о٫�o�}Z�\Q;]MBg2Zr�G� Y� {l��	�:�f�?���tj/�Ս��6Bj�!�`�(i3M�yx�,�G���V��H?Ә�%"Q�ܦfM� �L�Y}śT�!�`�(i3!�`�(i3G�&ց�*�p8�Iט��ō�Zm\�l��ì�A���V��H?Ә�%"Q�ܦfM� �'9�5���c(H޵D7W�:����p�A�ԍ'8����J�������"��<��y�@�v�&Sq�aj(��;����_��%$>_�n�To�[B���v�쟎��V��H?Ә�%"Q�ܦfM� �in5�҇�?�b��v݋N�����U-�pë��";Yy\'{w#/ B!�`�(i3޼QE1������m�(��k8һ��6ݕ��wp>�\�H��/Sg�Al�a�;�����9�Xy+�Mk��趵��1�F���������m�(��k8һ��6�D��)��	u�}�Q���GM�о٫��s�~�L�1{&��� )S���z;]MBg2Zr�G� Y� {l��	�g�yl��6T�T�D��ao.\C�kT���/T$ǩ����m�(��k8һ��6ݕ��wp>�\�H��/Sg�u-Y2�G�1{&��� �5掼�s��ݚ�Н�!�`�(i3K7͍��|��W&":!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�l~�1��n��+��o�JJ�tsq��T�G�'�q��;��y�-���2���澝ߚ���PC� �ˆ��*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��[��m�U����#3T��_�[g���pj������e�S�[�k]m��
ae���K��ʭ�!c����fx'v�ao.\C�k C�Mh�n �O`�Ag��ۭXX0���?V�#=uz��ɜڈ�KK?Ba���$_��v�z`��E�4ki��w�K��r�]�4�P�l��=5;���o�1g��U-�e'+]�{0C!�`�(i3!�`�(i3!�`�(i3AԢ�a\�g.��m6]c
j���%��g:���1nSpɃb6vJ�pZ� 4�F�Α��Bʏ,�:��O�?�I))����A�m�(�UVh�hP[�t��#��l��姹�xAQ�Y;x����$����7��=�S:t�L)��k]m��l��e b6vJ�pZ� 4�F�Α_)'!��r���U�4�8�v1a{J�j�f�AtT��_�[g�����,��WdM4@��_�U*��{��������
��\�H��/Sg�w��'o�GM��QО��i/R�c� }!�`��8
|�Kvb6vJ�pZ� 4�F�Α�v1a{J�j�f�At╔����̞��>��b��v݋N���������L+-�8���/����̜�I0���ԏ�.fOe	pۙE�����WdM4@��_�U*��Wc��V9a�Fc���M똡���iA'R�	s��]C�m�(��k8�4k_ł�k]m���E��Y� ,���� ��̆���M똡����o\�B/�u���a�x����r͖�1r����X�N�SF�vb6vJ�pZ�t���%�Q���� �^]�y܃fs�A���5��Q���� �^/s�1��p����;q�Zܑ��B$�䪜Q3N������2(wUF�|��: ��ao.\C�ktg����U��pqo�}9�-�_����NǨQ�~�^��>}�;�D#��2~��vNOgۈPM�r�]�4�P�l��=5;,��'ٕΖ�%����%2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�w�u��[�wbk�$�Z��Ջ`,9�H�W��`�z��Y��)h��{��Ķ�,�����F�!��cܦ���ҧ�v1a{J�)�3�� E!�`�(i3!�`�(i3�I����~u[��m�U�tV2�8�.�`��ai���Q��B%W����˩I4��欱���j���1#Y�p�� �VBD�!�Ĵ��ޯi��:��:̹��.�g3Z�7�4��~�U��{��0��L�r:h]��Ve.*�QN������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܨ$�`V1���cЉ�M�$@PJ+5*�轓�A1�J�����)����Ҿ���M���X���̜�I0���ԏ�.fOe	j�)6)-
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd�V3����C��z���Bf���a�x�G9�:Q����v�z`���pqo�}�;-�]�̓@?5�M%jWhC䨛��D)��C�V���3������G��������M���X�����9�;]MBg2Z�ܱ�Q3�!s!��xlJeYSWe^E1��b���t��w��X����xQ�1���~!�`�(i3!�`�(i3޼QE1���������M���XR����� ӫ/��mt����� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha3@��[/�������ܦR'cf���³5��*�7`����\Z��K�����5�O�%E#P����ҧ�v1a{J�"M�X�m�Z!�`�(i3!�`�(i3�I����~u}c��ko#���uT�.��=�F�@{2귑����|�kI��RhF�� ��*�C߇���t�k]m���E�i�m}66j�"Hs�@��C�,ԭ}3Y�Z��E��3?�d���&�Û=�������fo��ZpW4%"������k�I��RhF�䂔�R�D����M���XH {��u��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2����X�G[��7�癆cgQw�c4~Nr_�mS8<�n/�"����5=��)Q���nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��#�աl����aGl�97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��y���'j��ݚ�Н�i#\��u�vc�jj&��G�9m6�̟�1��"~6���aq��3=]��m�D��-����!�`�(i3px!��ia��T)�
���l�K�>�������Ra])n#���r����`
 ֢���̟�1dN�<@Iv��nt=:��:5A��pfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�ն'�U;|�� �R�SBJ���z`�3ޕ ���t�T��?E-h��`f���sd�G}%����3f闶P���`�3ޕ �7�癆cgQw�c4~Nr_�mS8<�n/�"����ZRR���dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ�0�p9zr��XƤ5_���"~6���aq��k�7� r��H�?�k ���50f
V��.ᬵy��f�'XĘ��L�F.	-�L��&PY~�y����o)�T*�c���-/a8!�`�(i3닓.�`�3E�g�������(ӈ���m�r����Ra])n#���r�����+��9,(ZRR���&���Ɗ3I5=��)Q�]� ���_�hbvk~�#x��	���"��]ap�~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�N(	I��^� �&����	cS�6�=P�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxִ/pJ��#��p,m��Q���M�"/���h|����6�o8:4�I���c�90��G��6�iI9�o«IX0F�M��uR3��%<�X�7�癆cgQw�c4~Nr_�mS8<�nQ'݀�=�Xy+�Mk���[��9�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�鞏̩jv�^������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��JFХ�B�9�4br���qP�V>t'�̗����S]�_�_��u��r��M�yx�,�G��i/R�c�'DV���b�z'hۉ)��d�7�q�՝� s�#���k$ �H�����4br���qP�V>t'�̗�����F��~1tSjv�!�`�(i3Q�>�H�((��"Jk�\p��j�������\�z�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxlP�6=��Nh�����x@�*�j��m�(��k8H {��u��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\75�e��4��X�G[��7�癆cgQw�c4~Nr_�mS8<�n(�6k�4dFn�H�~M�h��,���ANʂ��t�Ǌ���z
A��Φ�gz(AٸI))����A�m�(��2M�`�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�鞏̩jv�^������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��JFХ�B�9�4br���qP�V>t'�̗����S]�_�_��u��r��</Sn���̟�197��EN��~�{�B��R��� �hvT�+]�x}NI0���ԏ�.fOe	��;csj/�՝� s�#���k$ �H����p��j�����8"c��"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3��T��xW����˦G�m�(��k8��0�m���!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�Mm�(��k8��xh�j�W���5L5@�m�$R�nS�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2���j"�²O�i.����bs��2[�a��o���H�RtV�^G9�:Q����Z$�x$�֯� W97��EN�Q,�SGŹ�R���/�O��� ӫ/��m�A0`��A�2�����$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&r#o�]�ʄ�g�s���������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��;�uO��Bu����aGl��Z����pG�p�P�m������� h�ҩ�޼QE1��v1a{J����nFy� �����&��"]c�#y�>�)L�����/s=s�^�?��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxģ��_�ڑ��� en��`��n5��=�8�`Lv�RU��n;3ѫIX0F�MV�ҁGG%4vkz����`���φ��<�6�15���Dl=*�QN����r$ɓǃl[�Ƶ�1tSjv�޼QE1��v1a{J���Ꭓ�[��^E4+у��b�Bϱ��b��v݋N������M}Ĭ��ʡ.,�-��̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q��Y����(��U� P"G�wk��M똡��A�{�>�� ��
^�Mi~_�THN��R��bP�63Z�t�5ߧE4��Fr��j����bm&����T���Ꭓ�[�"�2�~�m�ek�}/�*��^��φ��<�6�@a� ��fFMqlg{y����i�q,?5qi��(.�j2��w�V�"xjzӝ���I(͂��-����N��r8!�k]m����DބiM�^E4+у��b�Bϱ��b��v݋N������M}Ĭ���՞)Ǭ�Q̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q��F��P�?�u�$�+AԢ�a\�]c
j���(y�.
جH�)��
���z#��#��Ě����E�i�m}6O�D mWN��ܐ�}��s����$c���Dx<�Θy9����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�޼QE1��v1a{J����nFy� �_Y��t��3
�v�v-}�	mp����/�כ�"]c�#y�>�)L�����/s=s�1�3���3
�v�v-}�	mp@?��jV�H�I�_Pg<���7�*w�ɝF�l�u�*Ha���J*�Rs�0�ǳ7��y.+�F�$-�S:t�L)��k]m����\�6�=�r��J*�Rs�08�b(��g]�6��;b#y�>�)L�^b٫
zܫ5u�q��	�����aq��p�Rdae�Qטg�u2]c
j���(y�.
جH�h��p\��"~6���aq����{M�jX Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������N��r8!�k]m��5L5@�m��i�*O����Qטg�u2�Tt$Ó6N�֤���n���6����?R����� ӫ/��m�A0`��A��7A�Ǩ�3
�v�v-}�	mpBR9ƭ�����fx'v�ao.\C�k�ף�D�~.8s�Z��N��r8!�k]m����\�6�EM?�ۄ�a�x�]c
j�����7�*w���Ǌ����fx'v�ao.\C�k�ף�D�~��pr����)x�?{���x.�Knq��!cI͸I))����A�m�(};l�-����׭�i�#�}��il��Rm�㭼�S}�S��S�C���+�%�t�*#y�>�)L�^b٫
z�.h��E��B\�H��/Sg޶��g�R6Ӹ�m ޶&�hbvk~�#x}���y���>��� ӫ/��m�A0`��A�;��ܞt�td���52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q����Z$�xQ�RY�##�� �~�^#y�>�)L�����/s=s��4�+��_��A5W��v�8:D�!�̞{��L]Eц~_�֤���n���6����?��ө%�Sg()��ikp���H���]c
j���4���TS3���/k���m���+)x�?{���<m�N=-�w���+ާ�����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3G9�:Q����Z$�x�vG��*Ha���J*�Rs�0K=X���d���fx'v�ao.\C�k�ף�D�~�Y�I���I�_Pg<���7�*w��D��q��� �~�^#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<���7�*w�ɝF�l�u�*Ha���J*�Rs�0��|�_�Y�j�W����΂o�����4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J����0;�����5u�q��	�����aq��ɪw�*=>@\�H��/Sg޶��d��5��f�C�7ª6��J�������ߧj@QEM?�ۄ��I�_Pg<�(y�.
جH��O��U
hPߺ0��A���ۖC�#dG訠�O`�Ag�v1a{J�Bz��s�V��m���+)x�?{����}9��|�G9�:Q��F��P�?��4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J�������ߧj@Q�_Y��t��3
�v�v-}�	mpl�!����_�n�To�[r��}k:�2Y�ا 2'l:}��Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc]�&P��	��I�_Pg<ˉJLg�2'�r�G� YF��6�!�`�(i3!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Y����G[�����a�x����r͖�k���$,�C�7ª6�{V�-_8���G�7W�:��G�z㤧{��B��+ H!�`�(i3!�`�(i39a�Fc���M똡���֤���n���6����?���$����;-�]�pR�$5iL�Pf8e���N��r8!)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��J�a$�Y �������G����1�E�AvY�5�h�B�c\��L̎C��fx'v�ao.\C�k�ף�D�~�Y�I�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��[�t��#��l��姹�C�`N���$@PJ+5zqiS�Q#y�>�)L�b�@_	��}Pz1Z�ݗ�"��I�����f�l��=5;R�ˊ	18kQ����&|���BY��l��=5;R�ˊ	18EYx��*��O`�Ag��ۭXX�|ʡi�����Fz�!�`�(i3!�`�(i3����&���0���y�هj�W�����ד*(�os}�&à�m�(��k8�*�0�mI0���ԏ�.fOe	m���h�����̜�I0���ԏ�.fOe	m���h��֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@�k̇���AEM?�ۄ��I�_Pg<ˉJLg�2'�r�G� Y�ҹnЭ:��#�@����ۭXX���E��O��j�W���bԽ�b��˔ �y=kg�������8�`Lv�RU���7xw���	�e��1{&��� �5掼�s��ݚ�Н�!�`�(i3]c
j��ʉJLg�2'�r�G� Y�)�?���I))����A�m�(};l�-��	}�<�Q"!�`�(i3�����9�Xy+�Mk��L

�F����8�`Lv�RU���7x�.9�?	��j�W���bԽ�b��˔ �y=kt��w��X<���H1���~!�`�(i3m��i�*��{V�-_8���G�7W�:��G�z㤧{����+c_�n�To�[r��}k:�>�hyȷ����wP?��i/R�c��;=~.�"�f!Hb�G����1�E�AvY�5�h�B�]�{���j�W���<�'��V�I�'��x!5�kz���[h�x�1W0�u]9�#�I���jVѭ@!�`�(i3 #��zG���{V�-_8���G�7W�:��G�z㤧{��B��+ H�ݓ�W���"r�DyA�S⏸[��t��7�M~G9�:Q����D����1�Q�
w�8D�t�%o�V\�Z�0��{V�-_8���G�7W�:��G�z㤧{��ԍ'8����J�����"�f!Hb�G����1�E�AvY�5�h�B�$5z&�D���ME�R�, �5��U���j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR���bn�u]9�#�I���jVѭ@!�`�(i3 #��zG���{V�-_8���G�7W�:��G�z㤧{�E2p��F4F�[��\	.���#�"r�DyA�S⏸[��t��7�M~G9�:Q����D����1�Q�
w�8D�t�%o�V\�Z�0��{V�-_8���G�7W�:��G�z㤧{��ԍ'8����J�����"�f!Hb�G����1�E�AvY�5�h�B�$5z&�D���ME�R�, �5��U���j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR���bn�������mo��jVѭ@!�`�(i3��dN���ub�z'hۉ)S���o޼QE1���Ꭓ�[��Yi䚠�5���u�L�!�`�(i3!�`�(i3!�`�(i3��c���鿉�X+�kQ��v1a{J���Ꭓ�[����$����;-�]�pR�$5iL�z#��#I	�����g[�s6{޴�i��)���!D������eW�d/=me�%b\%�I����~uI	�����g[�s6{޴�i��)�������T�\�H��/Sg޶��d��5��f�C�7ª6�)��%��+b�O~1��GM�о٫�S��wE\�!�`�(i3!�`�(i3�I����~u͘6��q���j�W���yͧT���E����ua�����\�ec[�U�b(l�rD��ЀUg]�6��;b�����5qo��o�����&Sq�aj(��;���Q�y�QF��fK�Ěk.�����GBz��s�V�r�G� Y� {l��	�m��ze��I))����A�m�(};l�-��o���n[�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q�K�\7}�W,��+G���*�1S�@:8S�C����0���y�هj�W����΂o���R��o�3��rD��ЀUR����� ӫ/��m�A0`��A�"��(ޅ���>��� ӫ/��m�A0`��A�,���$�n�M?��hS⏸[��א �k/ׇӭ��!�`�(i3!�`�(i3!�`�(i3����}>R� [�'a,�v1a{J��¸�k�Lpަ	<�%�;�ÇI���fx'v�ao.\C�k�ף�D�~���~�C9w��fx'v�ao.\C�k�ף�D�~h1��'�t�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��⒍~��Ĵ��ޯi��ŁO�(K���}�H[W2q�[�Kx�ʁQ7W�:���iޚuq6p��j����Q�9�|`ЉɁmwl��\�6��#P��Ѐ�5�h�B��ME�R�, m��
~�B�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\����oW���";Yy\'{w#/ B!�`�(i3޼QE1���Ꭓ�[��Yi䚠疛!wFii��{s��ֹ�Em��r�~ʁ���Mյ��#�@����ۭXX���E��O�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\L�}��鋿 ��
�Q�
w�8D�t�%o�V����������F>�w�γ~<�����6Bj�!�`�(i39<��`f�R(R�X���Ǹ���m�(��k8һ��6�R����� ӫ/��m�A0`��A�,���$�f��EJ,�G7```+�ֶ������]G��܎~:Q��z�˔ �y=k�2�u��܉�ӌ$/k�Bz��s�V�r�G� Y� {l��	�:�f�?���tj/�Ս��6Bj�!�`�(i3M�yx�,�G�����5qo��o�����&Sq�a��z#׊;w!�`�(i3!�`�(i3G�&ց�*�p8�Iט��ō�Zm\�l��ì�A�����5qo��o�����&Sq�ae:rmv�H�!�jT7|�`\%��u7W�:����p�A�ԍ'8����J����T"O5�`�7B��[�<?Ә�%"Q�ܦfM� �in5�҇�?����XzRL��MWX��DބiML�瞩w�j���@ΙN�[���-ل�{s��ֹ��!n)\HL�U���W�H�2^�/3!�`�(i3�0�9&،�R(R�X���Ǹ���m�(��k8һ��6��b��QM!Ϊu��U)�(*�O�q�@��i)&
�k�����oT`kz�)��%��+b�O~1��GM�о٫�o�}Z�\Q�R(R�X���Ǹ���m�(��k8һ��6�^?���I�^$D��Ҽ]G��܎~:Q��z�˔ �y=k�2�u���e�՝*U��eW�d/=4��b�Bz��s�V�r�G� Y� {l��	�g�yl��6����������F>�w�γ~<�����6Bj�!�`�(i3=��a���my$�N��o�/���;B����WN�Q���=�&�Φ�3h]��Ve.vrWB�i�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܧG%�MP3ö�3���Cw�Hm���9��N	{8G9�:Q��F��P�?\��R?��f�I))����A�m�(};l�-��Y��bq7h9��n� I�&|���BY��l��=5;R�ˊ	18�׼�^`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��I�_Pg<�(y�.
جH��O��U
h�07�;|''����˦G�͘6��q���j�W���yͧT���Ek�s���qa��;���=��i�uP=�z�}o*o���D)��ʱ�O�Ϸ(K���}Ǉj�W���yͧT���E��UH���4�����ˮ�N��G9�:Q��F��P�?��4�+��_碍�(H��(�K��k]m����DބiM�YG5`FFB���r����+C�ާ�����ݚ�Н�!�`�(i3!�`�(i3�I�_Pg<�(y�.
جH��O��U
h�07�;|''�)�?���I))����A�m�(};l�-��X;l_��Z2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq]�~��B�56e����bn3�qj]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7������B�56e��Y�p���]nA(�c���_G��Hb� h�ҩ�G��-�HG(�b�'Be���0��_�,\��݇��h	��F���L��b��v݋N������M}Ĭ��ʰ"���(���B����: ��ao.\C�k�ף�D�~��(��ᩁ��@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*�Va�ir���M��2"���&�^��v�8:?�'��ᦾ�;���8���U�._�nQ�rV��q�t7�v�]��1���U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^��@�z]��C�x!�H�k��^)(���27:����i�k�G/�����	^%�R��^�Mi~_�THN��R��bP�63Z�t�5ߧE4��Fr��j������B�56e���D����a�.m��K�+���w�?�H$~��	�����aq����>s�P�T����ym) �S���}�cЉ�M1y���TJ*�Rs�08�b(����Ph���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vck�ss:mo3G��-�HG(�b�'Be�i�}���$@PJ+5y*���� �S���}�cЉ�M�V�O�SFl�A���ۖ��S�<Ԣ������f�l��=5;R�ˊ	18kQ����&|���BY��l��=5;R�ˊ	18�׼�^`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcb��D�/�����	^%�R��aX��͟i8��m�q�/��v1a{J��U�Iv}տ�:
hbvk~�#x+[.Sk�NAG��-�HG(�b�'Be����\)Pߺ0��A���ۖ�w㌐g�߂.m��K�+���w�?�H$~��	�����aq��Ż%g�VƇ�m���Ar)���r����!�`�(i3!�`�(i3!�`�(i3��j�4��k]m���k�����A5W��v�8:C��4�I[��I))����A�m�(};l�-���j�	30�����Q��B%��>&ޝ�?1P��C&��b��Ɔ ����-˄�_-����dA�>�[E��1���~!�`�(i3!�`�(i3!�`�(i3-�E��%��v1a{J�a
�E��`���:�#�.��N�x%�M�RG�_`��z7{'#O�v1a{J�����ciA9*�"FP��� �mD��.1|��I�����V0�k]m��������fQ:b׻���3�v1a{J��bC�������N���� �VBD�!�Ĵ��ޯi�`͘�c�N&��H8|2�c�P�@��E�)�`L��%P��,���|�������[�i�*���1���"D���;�Ӏ�<qs��#�����M<E��'Z*)�?�R��n��h
:h����t�h��W+��W��v1a{J���&Y��V�Ԙ~q�9����t�T��?E-h��`f���sC>��Ӛ��S�J\7&���"�g72O!j���v�۲=�k2;�jmT�#bs��2[�a��o���H�RtV�^�G%�MP3�;ƹ��:i!�`�(i3��nF���<�W�.�P�	��
�Q�}9��?xs}�k�����|	�WIx����E2b�z'hۉ)��d�7�q�</Sn���k]m��D+_{6/ ���we��0�U+�qbp@�!�`�(i3[��m�U�H"҆>X� ��H�B�{_8�Y��=�}�Vݨ��}Dq�f��⒍~����v�z`��Ǖ��`���nF���<�W�.�P�	��
�Q�}���Mڷ��iA'R�	z�#,gB��3|v��Eb�z'hۉ)��d�7�q�Dw\����.m��TDZ��O$/ ���we��0�U+�qbp@�!�`�(i3�Ɔ ����;ƹ��:i����;q�{_8�Y��=�}�Vݨ��}Dq�f��N(	I��^��@K�]�!�`�(i3��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�G%�MP3�;ƹ��:i!�`�(i3���G��x��?�S��K�+���w�M�7��<�1�����\�H��/Sg�w��'oª���#oM��:<��j!�`�(i3�G%�MP3ö�3���!�`�(i3���G��x��?�S��}�k���ޗb�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J��湮��}6�/S� ����,��WdM4@��z(�ﳍ�f�_��S�>�!/�_�n�To�[
MQ9�F���"X��[�,�!���D!�`�(i3K�\7}�W,��+G��ܢN��_;��(���27:����7D!��%��g:���
A�%�q���F�dH�/�O��� ӫ/��m��M���	a(􆿳�3�m�
2]�!�`�(i3[��m�U/|w~S."����ʲ�P"G�wk�#�_wU|�1��v�z`넥^�?��F�dH�/�O��� ӫ/��m�A0`��Aw�zɝ8c��g��U-�e1�S������/��@���WdM4@��_�U*�u�$�+AԢ�a\�G�n봈2=��+G���*�1S�@:8M�7��<�1�����\�H��/Sg޶��j�}a�cf��"X��[�,�!���D!�`�(i3G��-�HG(�b�'Be��O����}ߟ�r�Q�C�x!�H��Yů�a��(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/���}Dq�f��G�dE�h�k]m��!�`�(i3g��c���b�'Be���I-�X!�`�(i3닓.�`�3BڴQ��J�a$�Y �Mn__��q��ڍ$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��'�al��p\ٿ�6�P)� &�]?�t�ϗ;��|B���?#�+Fz��Ԥ�Ԙ~q�9�C=2崝��tw�i�՗[�:X#x;2z��
�@h�5,Wlr�r%)cA��z>9�R��d���!i�6�5�p����M����-)O^��� �F��s]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M�v1a{J���&Y��V�scX{�X!,�'ž1�|�'����u��r��9��?xsTDZ��O$!�`�(i3x����E2b�z'hۉ)��d�7�q�`
 ֢���k]m���Ǖ��`�/ ���we��0�U+�qbp@�!�`�(i3[��m�U����L�F����;q�{_8�Y��=�}�Vݨ��}Dq�f��⒍~��Ĵ��ޯi�ʌ	���bS��nF���<�W�.�P�	��
�Q�}���Mڷ���o\�B/���2�>x����E2b�z'hۉ)��d�7�q�</Sn���k]m���E��Y�%��W#<e��0�U+�qbp@�!�`�(i3��j�4��k]m������;q�{_8�Y��=�}�Vݨ��}Dq�f�W����GTDZ��O$!�`�(i3��nF���<�W�.�P�	��
�Q�}����FYs96j��
!�`�(i3x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^9��?xsTDZ��O$!�`�(i3�i�<�~�y�j�q�7�AԢ�a\蟴���P`��ɠD(c!)��w�K��r�]�4�P�l��=5;���o�1g��U-�e1�S�������6���2[QvA�LO�>��
�I����~u�4br��
�uݟ�x��?�S��}�k���ޗb�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J��湮�ձ������r���IbW�P"G�wk�#�_wU|�1��v�z`넀r?&��AK��sC宸I))����A�m�(�QNȮ���k/��m#��}Dq�f����Mڷ��iA'R�	�yvc�]k�i�<�~�y�j�q�7�AԢ�a\�G�n봈2=��+G��܇�c.}M�$(���B����: ��ao.\C�kf��_@Z��T�\ �͆�v�9��</Sn���k]m��������fQ�qr�~�룺���aGl�k/E΋*U���7D!��l��姹�C�`N��䍬f�_��S�>�!/�_�n�To�[r��}k:�d4��f��a(􆿳�3�m�
2]�!�`�(i3[��m�U�H"҆>X�\2�~|G��YN
��)e
�����z%t��#-�v1a{J���!<�b�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p;�x'_|~� �S���}me":l�n�������r���IbW�G��-�HG(�b�'Bep�w�{�̞��>��b��v݋N������M}Ĭ���F`���G���`y����ݚ�Н���nސ�Ѵ����-VL!�`�(i3��DKY���k]m������W�!�`�(i3I8�ѐv2zigzA=v)����;q닓.�`�3��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�v1a{J���&Y��V�kcZ�Z�f��;_��8W�w��fD��e���WƂ�\���O�!2ɵ��w�o��'�R<l�K�T�}�̖˄��O��r��'������ܦR'cf���³5��*�7`����\Z��K��qb	��G��W+��W���fy����φ��<�6�@a� ��fFMqlgd�G}%����3fEa�F��x��A�Z����r$ɓǃl[�Ƶ�1tSjv�-�E��%�k�Vx3G�)P<�ܓ�Y�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&rG��Hb� h�ҩ�-�E��%�k�Vx3G��Mn__���ͥ
ݐ����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�Ea�F��x�j���NC�V��	��y���B��у#Y�wP-�H1�m��d�7�T
u�/%F���J���rG[Pt��H {��u��]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�Ɔ ���Ve��˅�E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/8"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3�p�8H���v1a{J�ikl(rco��(`��ү/�O'�=�CyQ�/Ap�H�RtV�^�G�dE�h�k]m��Cw�Hm���Ɔ ���Ve��˅��ԝy'��Ra])n#���r�����G�dE�h�k]m��Cw�Hm��K7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6����:��1=���N�KRoY����#�`18vP�� ���Jx�y�Zgl�fb�l����t�h��W+��W��Ɔ �������4�Ք�R'cf���³5����U��+�Xa�H(�˕�Eo(d�J��:�����nސ�ѽv1a{J�k�Vx3G�������S�CП�HN��R��?�d���&�N��	�Ȓ����vm��.�g3Zdj�t��a"�6�m��C������06S��^����$����2�"�1	�<����ߙq�|�����Z��㽕���䕠�s�����혅vº�w�⽒���M���o�G�m�?$��̼�K���Z��㽕���䕽v1a{J�k�Vx3G�(���27:��`.��5��C�)���t�Z����S�CП�R��X鷴QW�w��fD�Ɔ ������&e��c���L}���1LdO�{PH�b_�C���#<x=aUh��������-VL��y���[��,_���p���,@��a��NYs�����4$�[�l��~��R��ƿ;W ��.���:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�d�@���GE�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����4br������Ľ����Չxv��Օ��qvdЧ^{�j����'�����Z>ؼ��XyH�RtV�^�G:w�䖬n���~�����q�ZLN�	��MdGN���!�`�(i36�ZV	�	ҙ���˦G��d�@���G6 y2��R�՝� s�#���k$ �>=���#䖬n��؂�nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j �_�ȇL�X Hz��0�Jw��3�+=�4o���+��+}�K=���e���Օ��qvdЧ^{�jM|�"D5�O�%E#P��=m緒1d�;q3�)�U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩΟ/��mS%y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�	�)��&ghRV��R���P�|T����{7�H����8���O�υ���YN
��)e#j�o����:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�I��� g�����Օ��qvdЧ^{�jMdGN���!�`�(i3%Q�[�J����˦G��4br��6 y2��R�՝� s�#���k$ �B�'��a����aGl���nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN!�`�(i3]���-_!Q���ŴIh�5,Wlr�r%)cA/�r�]/2�ݚ�Н��ߎ ��E�VTҝD!u���o���F������}Dq�f��	��x��ݚ�Н��ߎ ��E�VTҝD!u��nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�k��{`.~��No�ߏ��T�4(���;��|BJ�U�� �X�G[�wE�=p���4br����3v�qh�5,Wlr�r%)cAQ17�b�����d���!i�/��mS%rƂ�o��+h� ��6j�"HsP�����X�G[�OL��qt�Z���#���2=��h��IX0F�MV�ҁGG%4vkz���յ[+8��r$ɓǃl[�Ƶ�1tSjv�>F��3��mlr�{��|e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3�}�P6@��e��>��Օ��qvdЧ^{�j@��C2K�ǽ$�!b����#�GWW�<om���濫�L��� h�ҩ��H�������M��2��22= ��v�8:?�'����-����!�`�(i3}�1�Hz8�ZF�*�Gx�����}Dq�f��	��x��ݚ�Н� ��4E|���Bf����{_8�Y��=�}�Vݨ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}Ĉ7NU�.j��u�Nb�BHn̐2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�S*�"�=3�Ҥ�P�X��������3R��kѶ���� ��&��h�?i�H��}��?<����G&�;���� ����}p閭3u��N�,?��΃���]�X�ֻla�oZx�i�xx�j�甯�[���pФq�Ǒ)''��m�9X��W��� �_%B71Ձ"�Ĭt�'�ǅ@s�-6��P�%Ae!�`�(i3<�6�Q=������Kd���{J��&�)HVi�pz��AY���Z�@���v��d�-td'�I1L�S���%�4/�p_�g�P���V�Wb<�..�4���ho7L��2�"�G�p�Pڹ��/^�w?�d���&�N-Y&yo�q��=m緒X�X�pF�{_8�Y��=�}�Vݨ�ʥ��F��|����"�`Ec'�\Y-φ��<�6�@a� ��fFMqlgd�G}%����3f���K��M�ZP�����V��)�)��H����Qw�c4~Nr_�mS8<�n�ݚ�Н�ʬw�S���q9+t�}�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv������$ɔ9Q<ϯXr&ߜ����>05H~
�:qEp�;�P�t�5fĉ>99��A0ok�׹�x+��IhШ��+���Al+�H�A[�á��'G�+p�Dʾ��6�o8:4�I���c�90B3v�A��{y����i�q,?5q�+�#4��F��8M�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�2VP��Ѣ2����L��my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�<�i�������M;C��!��iKk�������J*�Rs�08�b(����<��#�!�`�(i3�j���%�|�;�ƇT��J��sr�l�ԝy'�fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx'X���5����'G�+p�9���?�(�JZ�Vk�;��|B��loXBȱg�S>X;Z�˯��R����e���Wƍ ٻ�l���M���R��ӟ-���4�&����Z����`	p�=�3Yj>�B�R���$]'\gWg��	�Z�kfc&�2���� ��b�FP&�r�@|�TԼ�\�v��_�R�GO.C�U��B��-����A�;�����\�5ｵ����;�jmT�#bs��2[�a��o���H�RtV�^*�9��.����N�eM�#��}Dq�f���NƥNoz��KUq՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r���'��o�u:��_x���O����]�!��	Ǹ�y85��8��,	iL�*dgN;ۍ����$9���Z��o�^��D���:5A��p��(1l�jG���Z��o�h�G KH�F;p�	%Ɏ�Bi!�`�(i3�ݚ�Н�-��)'���N�R���Va�irl�
@\�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н���������ۥ�Y�m���NM���!�`�(i3-6���[��<�p��Ar�8w�B
�:qEp�gdq�_x����Yzw��(4G��>��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3>�Q�c6���*(H=�ƍ2���l�!�`�(i35���u�L����˟y!�`�(i31���~!�`�(i3ʬw�S��ht��p���j��8�u��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��}�6�nq�Z�@���v�_{ޣ��$7������φ��<�6�@a� ��fFMqlgd�G}%����3f闶P���`�3ޕ �|#HK��A(�c���_G��Hb� h�ҩ�EOJ�uxm�7d��2�4.K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/8�@�����2
xH��!�`�(i3CT�MZ�\�XƤ5_��,\���*s-�e�2>J*�Rs�08�b(����T�\yb�����Z>��A�$�|��'T���+�L�F.0D�	�I���_
�u�����|�G�p�P�C������H8Џ�Ӿ���yi�1tSjv��wӨj]h��J��sr�lv{��lw	!ݞX�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�Mn5�b	���J��sr�laT��3G?�d���&����*�����E��h���O�Zj�������1φ��<�6�@a� ��fFMqlg{y����i�q,?5q���D5P��wFlE� ��'ž1�|�'����u��r��i��H�p��ic)�̩ƍ2���l�*�9��.�ԫ�&Np;qƍ2���l�����g�Z��3��a���!@�f")u��r��܌;���'����u��r���=�$���Ly���Cʬw�S��ڏ"/��z�>�Q�c6��?��!�6ʬw�S����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ���D5P�����+C�!-T��T�^���h�.k�mb�&��ƭ������xO��̋{b62�tstF�!��cܤ|�)՜�45�[՚1Dq��P�<
[�л���7Cw�Hm�̶^�+3���e]�#�?4�s_o#�{�U��)���Y;e�iK!���d.�% ��\:Fa�7�����~�L�D����C#/<���q�r$ɓǃl[�Ƶ�1tSjv�����,<��c�!{p85E�g�������(ӈ���m�r��������x���^a�nu4Bޗ��jw�	��C#/<���q�
�t��T&���LQ�/81tSjv�k��u������}�Fe��1�:��g�XW-#��=���;�P�t�5:Ha��VK�;�P�t�5E�xa�/ݺφ��<�6�2VP��Ѣ� (<ݐ�k-|���vG����и;2z��
�@h�5,Wlr�r%)cA��z>9�R��d���!i�%ؙ,{F�}�1U��VP��t�i?�i2�.[W�w��fD|�O�E/�Ĳ�=�Z���^��[�n�2o� #�����M<E��'Z*)�?�R��n��h
:h����t�h��W+��W���ŊPTWo9���gѸ-���֫IX0F�MV�ҁGG`5:�����+�^n=\f�5>����Db^<�..�4��<qs���|#HK��A(�c���_G��Hb� h�ҩκ%ؙ,{F��#QSU:�����|e"�O)�b�c�!{p85E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н��%ؙ,{F���\D�E��hW��ڬ!�,���6+�<�6�Q=5����.������w�h�8Vb5����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī��K��M�ZP�����Fz��Ԥ���엝�����L}�]���4x;΂��m9Ϲ@��2��w���.�
���t�T��?E-h��`f���sC>��Ӛ��S�J\7�p���"Z�v��!;�jmT�#bs��2[�a��o���H�RtV�^��~Щ�%��v��՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!�Bt�wz3��0��I8�ѐv2�_Y�d��o��b�Bϱ��z�
����{�g=_[�7����닓.�`�39����6��ݚ�Н��L&�Ǟ��W�VL��׬��P�|T���nT����
y���^��D��G��q"Y��;����rx�pj�d!�`�(i3��Q7lY��u�M�Һ����1)uם�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j0C.�>��VaT��3G?�d���&�<��vQ�zi��Hy�GE��R���H"X�0��n���l�IX0F�MV�ҁGG%4vkz����`���φ��<�6�Q١Ӿ�$	��1�h\���F�`yx�>�+X�M?��y�Bz�;{/�>��]#�y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�Y�)�}��EXs70��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��a�F�������Y���D��3��b�]결���:$�O���jF�ཕu�_�mS8<�n�ݚ�Н� �#0xg�`�I��Wz}�ἱc��-).^QQ�b��~$�
�:qEp�;�P�t�5����l��~��?�kv��.V��:��������kB�����X!o%�ſ����O?����<�5�>�?�R��n�K��$�<ۧ�: ��ao.\C�kFGˤ]u���:����
�ݚ�Н��>���Dl����|�b�и|��?���a{�w�!]��̍��}Dq�f������!�`�(i3oj�+p�K�J�iN�SE�g�������(ӈ���m�r����fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�Ӫ��*$���A����ƃ�Y���D��3��b��-��|^a�����Q١Ӿ�$�XƤ5_��,\���1�Hs�k���*��'���9���T�Q١Ӿ�$w���	�e���0��Qܓ'{w#/ B!�`�(i3!�`�(i3$ʩ�})��W��CX-+;X���X��ͷ(�-��]a;����D厺��+�XƤ5_��,\���q���7?�R��nI4�p� ^�b��v݋N�����AS�$�[���G��f#��O?���#j�o������6Bj�!�`�(i3!�`�(i3�����z!J��/٣��q8h��^�Q[M��P��#��s�'	�?��[��羹�He�-�c��R:k�ڛ���Ο]_Z鎬�����	�7 �#�E ���� ��M�#зq8�Ј'���Xw�P���w��a�e56<�5{ΖM+����+�J���q���U��D�U�2Y��i�p��+�FJ�9��V��Q]� _ό���.�@?d�s�8KFmғO�4}`L����D:�n`5�fK�\w��0]\o�LCd�|�w��DK����$���7s�9���o>��l%i�-}�
�?�v�-���w:���z�Ji��d�٣��c�A�L'Qī�*pY�M�l��S�J*�Rs�08�b(������l__��E� )�&��"X��[��Q[R�7�$��Xo��� ���Lk�Bgt�#P4];ˍH��M��=�&&ĕ^$&�	�s�{܇����O�յ[+8�a�)��Ƃ~6T���Q�x1�~g_�,\ަ�It��+g[�Zt%��m&<>��%��JU�a�(�n����62�tϛA^��'T���+M�Mb�:u�w�vG�q�:�&����#|�1�0j��*������Э~���V��2
L.�X;p`��3
�v�v-}�	mp,��_А#�<om���'$W$�X�t����}�(�
4��c��^�
E����d���m l�o�&�C�/w�x�P���E�`JcU!�`�(i3XO����0¤լq��/,���9^-��X�0���X�q!�`�(i3���)�>�)x�?{���x.�Knq���;W��ZLN�	��f�?ǉ�=@�#=���ix���!�`�(i3��ԫrI�C�i�4��v�(��.��dLG���6!�`�(i3���K�7��1۳ఋ�ݚ�Н���*dy�ZB\w��B���!�`�(i3�)ύ^��R�^Ƒ��f�?ǉ�=s���eZ�c]��E���!�`�(i3Q)��Zl�z��SR:g()��ikp���H������7Pr��ġ��,�a��OY�P�CQ��Bރ;�{��C�{����K�7��C4%̈́�(�y�|����x��~iM5/�S3 <�X;p`�M���ʄ?�k�V�?egE�@��i!�`�(i3-��,%>ʴ����қDO,\ͨ܉p����O,8�ݚ�Н�7�N�-��#l'U:�g[q�vG+|�<竷b��"&�_~�:N�4�0 L?�p���@Z,�ttT��Q�#<4^�>N0Θ��ݚ�Н��0V32;5�-�����4)cq�vG+|�<?V��j�cc����L�{��%ў׫>V��2GɎ�#���?\a��4�czZ��������[�D���~�ߗ���@Tvs�!�`�(i3�$�~c/�R��ŭ�.
�:qEp0���Y$���/ӳxW8�8J�|9 �P���R�A��4�h���!U�020�$�~c/�*���J= �P���R�^=^���3!�`�(i37�_M���{�� ��YOZ@��5�h�ʪ%��18�$��`��UB�L5wG�!�`�(i3��2]��ٱ�R:k�ڛԀlY�{:fh�3�w�	�|�s�Õ�M�<���{L,8ԀlY�q-�~_@!�`�(i3�[�H���,޷��u�2�1�9~F�r�t��b���չ�Ad���Ô�b��N�[\�i�]���B��E, �c��ΞOߙYĸ-�4:� �
�	(��7��F�dHw(��ES���v�8:ۛ@W:���#���FӪ�c�g<�j"Xt�F�)��#L����@� ��X�u�%h�K��(�%�z��I��s�*2��3��Wғ��7��&���oC���T8e�i�������ᳮ�T���t�T��?E-h��`f���sC>��Ӛ��S�J\7�p���"Z�v��!;�jmT�#bs��2[�a��o���H�RtV�^��~Щ�%��v��՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�$XR�QܛOcOZail������&G!�`�(i3��Q7lY��u�M�Һ���BO#LB�q#a�_�̞��>��3
�v�v-}�	mp,��_А#�<om�����M��2;!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j�p���"��NwK�"�Q=C&pm" <{>w�\�S�-D�I��L�@��8Q	��+���XƤ5_�J�	�LÆ���#��k���Ϊ�iIn���I_�1����!�`�(i3��7I���aT��3G?�d���&��J�p�k���\�#�k��m6[��!N�'�y�G