// Swept Source Optical Coherence Tomography acquisition system
// 
//==============================================================================
// Copyright (C) 2011 LIOM Laboratoire d'Imagerie Optique et Mol�culaire
//                    �cole Polytechnique de Montr�al
// Edgar Guevara, Maxime Abran
// 2011/08/18
//==============================================================================
//  This code is generated by Terasic System Builder
//==============================================================================
`include "my_incl.v"			// Verilog include file

module DE4_DDR2(

	//////// CLOCK //////////
	GCLKIN,
	GCLKOUT_FPGA,
	OSC_50_BANK2,
	OSC_50_BANK3,
	OSC_50_BANK4,
	OSC_50_BANK5,
	OSC_50_BANK6,
	OSC_50_BANK7,
	PLL_CLKIN_p,

	//////// LED x 8 //////////
	LED,

	//////// BUTTON x 4 //////////
	BUTTON,
	CPU_RESET_n,
	EXT_IO,
	
	//////// DIP SWITCH x 8 //////////
	SW,

	//////// SLIDE SWITCH x 4 //////////
	SLIDE_SW,

	//////// SEG7 //////////
	SEG0_D,
	SEG0_DP,
	SEG1_D,
	SEG1_DP,

	//////// Temperature //////////
	TEMP_INT_n,
	TEMP_SMCLK,
	TEMP_SMDAT,

	//////// Current //////////
	CSENSE_ADC_FO,
	CSENSE_CS_n,
	CSENSE_SCK,
	CSENSE_SDI,
	CSENSE_SDO,

	//////// Fan //////////
	FAN_CTRL,

	//////// EEPROM //////////
	EEP_SCL,
	EEP_SDA,

	//////// SDCARD //////////
	SD_CLK,
	SD_CMD,
	SD_DAT,
	SD_WP_n,

	//////// RS232 //////////
	UART_CTS,
	UART_RTS,
	UART_RXD,
	UART_TXD,

	//////// Ethernet x 4 //////////
	ETH_INT_n,
	ETH_MDC,
	ETH_MDIO,
	ETH_RST_n,
	ETH_RX_p,
	ETH_TX_p,

	//////// Flash and SRAM Address/Data Share Bus //////////
	FSM_A,
	FSM_D,

	//////// Flash Control //////////
	FLASH_ADV_n,
	FLASH_CE_n,
	FLASH_CLK,
	FLASH_OE_n,
	FLASH_RESET_n,
	FLASH_RYBY_n,
	FLASH_WE_n,

	//////// SSRAM Control //////////
	SSRAM_ADV,
	SSRAM_BWA_n,
	SSRAM_BWB_n,
	SSRAM_CE_n,
	SSRAM_CKE_n,
	SSRAM_CLK,
	SSRAM_OE_n,
	SSRAM_WE_n, 

	//////////// HSMC-B, HSMC-B connect to DCC //////////
	// Data Conversion Card
	AD_SCLK,
	AD_SDIO,
	ADA_D,
	ADA_DCO,
	ADA_OE,
	ADA_OR,
	ADA_SPI_CS,
	ADB_D,
	ADB_DCO,
	ADB_OE,
	ADB_OR,
	ADB_SPI_CS,
	AIC_BCLK,
	AIC_DIN,
	AIC_DOUT,
	AIC_LRCIN,
	AIC_LRCOUT,
	AIC_SPI_CS,
	AIC_XCLK,
	CLKIN1,
	CLKOUT0,
	DA,
	DB,
	FPGA_CLK_A_N,
	FPGA_CLK_A_P,
	FPGA_CLK_B_N,
	FPGA_CLK_B_P,
	J1_152,
	XT_IN_N,
	XT_IN_P,

	//////////// HSMC I2C //////////
	HSMC_SCL,
	HSMC_SDA,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	GPIO,

`ifndef USE_DDR2_DIMM2
	//////// DDR2 SODIMM //////////
	M1_DDR2_addr,
	M1_DDR2_ba,
	M1_DDR2_cas_n,
	M1_DDR2_cke,
	M1_DDR2_clk,
	M1_DDR2_clk_n,
	M1_DDR2_cs_n,
	M1_DDR2_dm,
	M1_DDR2_dq,
	M1_DDR2_dqs,
	M1_DDR2_dqsn,
	M1_DDR2_odt,
	M1_DDR2_ras_n,
	M1_DDR2_SA,
	M1_DDR2_SCL,
	M1_DDR2_SDA,
	M1_DDR2_we_n

`else
	//////// DDR2 SODIMM //////////

	M2_DDR2_addr,
	M2_DDR2_ba,
	M2_DDR2_cas_n,
	M2_DDR2_cke,
	M2_DDR2_clk,
	M2_DDR2_clk_n,
	M2_DDR2_cs_n,
	M2_DDR2_dm,
	M2_DDR2_dq,
	M2_DDR2_dqs,
	M2_DDR2_dqsn,
	M2_DDR2_odt,
	M2_DDR2_ras_n,
	M2_DDR2_SA,
	M2_DDR2_SCL,
	M2_DDR2_SDA,
	M2_DDR2_we_n 
`endif	//USE_DDR2_DIMM2
);

//==============================================================================
//  PARAMETER declarations
//==============================================================================


//==============================================================================
//  PORT declarations
//==============================================================================

//////////// CLOCK //////////
input		          		GCLKIN;
output		          		GCLKOUT_FPGA;
input		          		OSC_50_BANK2;
input		          		OSC_50_BANK3;
input		          		OSC_50_BANK4;
input		          		OSC_50_BANK5;
input		          		OSC_50_BANK6;
input		          		OSC_50_BANK7;
input		          		PLL_CLKIN_p;

//////////// LED x 8 //////////
output		     [7:0]		LED;

//////////// BUTTON x 4 //////////
input		     [3:0]		BUTTON;
input		          		CPU_RESET_n;
inout		          		EXT_IO;

//////////// DIP SWITCH x 8 //////////
input		     [7:0]		SW;

//////////// SLIDE SWITCH x 4 //////////
input		     [3:0]		SLIDE_SW;

//////////// SEG7 //////////
output		     [6:0]		SEG0_D;
output		          		SEG0_DP;
output		     [6:0]		SEG1_D;
output		          		SEG1_DP;

//////////// Temperature //////////
input		          		TEMP_INT_n;
output		          		TEMP_SMCLK;
inout		          		TEMP_SMDAT;

//////////// Current //////////
output		          		CSENSE_ADC_FO;
output		     [1:0]		CSENSE_CS_n;
output		          		CSENSE_SCK;
output		          		CSENSE_SDI;
input		          		CSENSE_SDO;

//////////// Fan //////////
output		          		FAN_CTRL;

//////////// EEPROM //////////
output		          		EEP_SCL;
inout		          		EEP_SDA;

//////////// SDCARD //////////
output		          		SD_CLK;
inout		          		SD_CMD;
inout		     [3:0]		SD_DAT;
input		          		SD_WP_n;

//////////// RS232 //////////
output		          		UART_CTS;
input		          		UART_RTS;
input		          		UART_RXD;
output		          		UART_TXD;

//////////// Ethernet x 4 //////////
input		     [3:0]		ETH_INT_n;
output		     [3:0]		ETH_MDC;
inout		     [3:0]		ETH_MDIO;
output		          		ETH_RST_n;
//input		     [3:0]		ETH_RX_p;
//output		     [3:0]		ETH_TX_p;

//////////// Flash and SRAM Address/Data Share Bus //////////
output		    [25:0]		FSM_A;
inout		    [15:0]		FSM_D;

//////////// Flash Control //////////
output		          		FLASH_ADV_n;
output		          		FLASH_CE_n;
output		          		FLASH_CLK;
output		          		FLASH_OE_n;
output		          		FLASH_RESET_n;
input		          		FLASH_RYBY_n;
output		          		FLASH_WE_n;

//////////// SSRAM Control //////////
output		          		SSRAM_ADV;
output		          		SSRAM_BWA_n;
output		          		SSRAM_BWB_n;
output		          		SSRAM_CE_n;
output		          		SSRAM_CKE_n;
output		          		SSRAM_CLK;
output		          		SSRAM_OE_n;
output		          		SSRAM_WE_n;

//////////// HSMC-B, HSMC-B connect to DCC //////////
// Data Conversion Card
inout		          		AD_SCLK;
inout		          		AD_SDIO;
input		    [13:0]		ADA_D;
input		          		ADA_DCO;
output		          		ADA_OE;
input		          		ADA_OR;
output		          		ADA_SPI_CS;
input		    [13:0]		ADB_D;
input		          		ADB_DCO;
output		          		ADB_OE;
input		          		ADB_OR;
output		          		ADB_SPI_CS;
inout		          		AIC_BCLK;
output		          		AIC_DIN;
input		          		AIC_DOUT;
inout		          		AIC_LRCIN;
inout		          		AIC_LRCOUT;
output		          		AIC_SPI_CS;
output		          		AIC_XCLK;
input		          		CLKIN1;
output		          		CLKOUT0;
output		    [13:0]		DA;
output		    [13:0]		DB;
inout		          		FPGA_CLK_A_N;
inout		          		FPGA_CLK_A_P;
inout		          		FPGA_CLK_B_N;
inout		          		FPGA_CLK_B_P;
inout		          		J1_152;
input		          		XT_IN_N;
input		          		XT_IN_P;

//////////// HSMC I2C //////////
output		          		HSMC_SCL;
inout		          		HSMC_SDA;
	
//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
inout		    [35:0]		GPIO;

`ifndef USE_DDR2_DIMM2
//////////// DDR2 SODIMM //////////
output		    [15:0]		M1_DDR2_addr;
output		     [2:0]		M1_DDR2_ba;
output		          		M1_DDR2_cas_n;
output		     [1:0]		M1_DDR2_cke;
inout		     [1:0]		M1_DDR2_clk;
inout		     [1:0]		M1_DDR2_clk_n;
output		     [1:0]		M1_DDR2_cs_n;
output		     [7:0]		M1_DDR2_dm;
inout		    [63:0]		M1_DDR2_dq;
inout		     [7:0]		M1_DDR2_dqs;
inout		     [7:0]		M1_DDR2_dqsn;
output		     [1:0]		M1_DDR2_odt;
output		          		M1_DDR2_ras_n;
output		     [1:0]		M1_DDR2_SA;
output		          		M1_DDR2_SCL;
inout		          		M1_DDR2_SDA;
output		          		M1_DDR2_we_n;

`else
//////////// DDR2 SODIMM //////////
output		    [15:0]		M2_DDR2_addr;
output		     [2:0]		M2_DDR2_ba;
output		          		M2_DDR2_cas_n;
output		     [1:0]		M2_DDR2_cke;
inout		     [1:0]		M2_DDR2_clk;
inout		     [1:0]		M2_DDR2_clk_n;
output		     [1:0]		M2_DDR2_cs_n;
output		     [7:0]		M2_DDR2_dm;
inout		    [63:0]		M2_DDR2_dq;
inout		     [7:0]		M2_DDR2_dqs;
inout		     [7:0]		M2_DDR2_dqsn;
output		     [1:0]		M2_DDR2_odt;
output		          		M2_DDR2_ras_n;
output		     [1:0]		M2_DDR2_SA;
output		          		M2_DDR2_SCL;
inout		          		M2_DDR2_SDA;
output		          		M2_DDR2_we_n;

`endif //`ifndef USE_DDR2_DIMM2

//==============================================================================
//  REG/WIRE declarations
//==============================================================================

//// Global signals
wire 						reset_n;

//// Master template
wire						control_done_read;
wire			[31:0]		user_buffer_data_read;
wire						user_data_available;
wire			[29:0]		address_last_complete_read;
wire						control_go_read;
wire			[29:0]		control_read_base;
wire			[29:0]		control_read_length;
wire						user_read_buffer;
wire						reading_done;
wire			[31:0]		debug_read;
wire			[2:0]		error_data;
	
wire						control_done_write;
wire			[31:0]		user_buffer_data_write;
wire						user_buffer_full;
wire			[29:0]		address_last_complete_write;
wire						control_go_write;
wire			[29:0]		control_write_base;
wire			[29:0]		control_write_length;
wire						user_write_buffer;
wire						writing_done;
wire			[31:0]		debug_write;
wire						error_full;

// DDR2 200 MHz clock out
wire						ddr2_phy_clk_out;

// Power on reset
//wire						reset_power_on;

//// Ethernet
wire						enet_mdc;
wire						enet_mdio_in;
wire						enet_mdio_oen;
wire						enet_mdio_out;
wire						enet_refclk_125MHz;

wire						lvds_rxp;
wire						lvds_txp;

// A-line of 1170 Elements, each 14 bits wide
reg  		[13:0]			A_line_array	[0:`NSAMPLES-1];
wire		[13:0]			A_line; 

// 50 kHz A-line trigger
wire						sweepTrigger;
// 50 kHz A-line trigger enabled by LabView
wire						trigger50kHz;

// Position of the ADC sample in the RAM
wire		[10:0]			read_RAM_address;
wire		[10:0]			write_RAM_address;

// Data from RAM
wire		[13:0]			RAMdata;

// MSB to write dual buffer RAM
wire						dualMSB_write;


// Acquiring 1170 samples
wire						acq_busy;

// Acquisition of one A-line done
wire						acq_done;

// Reading RAM 
wire						read_RAM_busy;

// PWM for Fan and LED
wire		[7:0]			clk_div_out_sig;

// Receive signal from LabView to record data to DDR2
wire						enableRecording;

// sinus wave signal
wire		[13:0]			raw_sine;
// output to DAC A
reg			[13:0]			o_sine;

//==============================================================================
//  External PLL Configuration ==========================================
//==============================================================================

//  Signal declarations
wire 		[3:0] 			clk1_set_wr, clk2_set_wr, clk3_set_wr;
wire         				conf_ready;
wire         				counter_max;
wire  		[7:0]  			counter_inc;
reg   		[7:0]  			auto_set_counter;
reg          				conf_wr;

//  Structural coding
assign clk1_set_wr 			= 4'd1; //Disable
assign clk2_set_wr 			= 4'd1; //Disable
assign clk3_set_wr 			= 4'd7; //156.25 MHZ

assign counter_max 			= &auto_set_counter;
assign counter_inc 			= auto_set_counter + 1'b1;

always @(posedge OSC_50_BANK3 or negedge reset_n)
	if(!reset_n)
	begin
		auto_set_counter <= 0;
		conf_wr <= 0;
	end 
	else if (counter_max)
		conf_wr <= 1;
	else
		auto_set_counter <= counter_inc;


ext_pll_ctrl ext_pll_ctrl_Inst (
	.osc_50(OSC_50_BANK3), //50MHZ
	.rstn(reset_n),

	// device 1 (HSMA_REFCLK)
	.clk1_set_wr(clk1_set_wr),
	.clk1_set_rd(),

	// device 2 (HSMB_REFCLK)
	.clk2_set_wr(clk2_set_wr),
	.clk2_set_rd(),

	// device 3 (PLL_CLKIN/SATA_REFCLK)
	.clk3_set_wr(clk3_set_wr),
	.clk3_set_rd(),

	// setting trigger
	.conf_wr(conf_wr), // 1T 50MHz 
	.conf_rd(), // 1T 50MHz

	// status 
	.conf_ready(conf_ready),

	// 2-wire interface 
	.max_sclk(MAX_I2C_SCLK),
	.max_sdat(MAX_I2C_SDAT)
	);

//==============================================================================
//  End of External PLL Configuration ==========================================
//==============================================================================

//==============================================================================
//  Structural coding
//==============================================================================

//// Global signals
assign reset_n 				= CPU_RESET_n;

//// Ethernet
assign	ETH_RST_n			= enet_reset_n;

`ifdef NET0
input		     [0:0]		ETH_RX_p;
output		     [0:0]		ETH_TX_p;
assign	lvds_rxp			= ETH_RX_p[0];
assign	ETH_TX_p[0]			= lvds_txp;
assign	enet_mdio_in		= ETH_MDIO[0];
assign	ETH_MDIO[0]			= !enet_mdio_oen ? enet_mdio_out : 1'bz;
assign	ETH_MDC[0]			= enet_mdc;

`elsif NET1
input		     [1:1]		ETH_RX_p;
output		     [1:1]		ETH_TX_p;
assign	lvds_rxp			= ETH_RX_p[1];
assign	ETH_TX_p[1]			= lvds_txp;
assign	enet_mdio_in		= ETH_MDIO[1];
assign	ETH_MDIO[1]			= !enet_mdio_oen ? enet_mdio_out : 1'bz;
assign	ETH_MDC[1]			= enet_mdc;

`elsif NET2
input		     [2:2]		ETH_RX_p;
output		     [2:2]		ETH_TX_p;
assign	lvds_rxp			= ETH_RX_p[2];
assign	ETH_TX_p[2]			= lvds_txp;
assign	enet_mdio_in		= ETH_MDIO[2];
assign	ETH_MDIO[2]			= !enet_mdio_oen ? enet_mdio_out : 1'bz;
assign	ETH_MDC[2]			= enet_mdc;

`elsif NET3
input		     [3:3]		ETH_RX_p;
output		     [3:3]		ETH_TX_p;
assign	lvds_rxp			= ETH_RX_p[3];
assign	ETH_TX_p[3]			= lvds_txp;
assign	enet_mdio_in		= ETH_MDIO[3];
assign	ETH_MDIO[3]			= !enet_mdio_oen ? enet_mdio_out : 1'bz;
assign	ETH_MDC[3]			= enet_mdc;

`endif

//// FLASH and SSRAM share bus
assign	FLASH_ADV_n			= 1'b0;				// not used
assign	FLASH_CLK			= 1'b0;				// not used
assign	FLASH_RESET_n		= global_reset_n;
//// SSRAM

//==============================================================================
// assign for ADC control signal
//==============================================================================
assign	AD_SCLK				= 1'b0;				// (DFS)Data Format Select = binary (0)
assign	AD_SDIO				= 1'b1;				// (DCS)Duty Cycle Stabilizer ON
assign	ADA_OE				= 1'b0;				// enable ADA output (active LOW)
assign	ADA_SPI_CS			= 1'b1;				// disable serial port interface A
assign	ADB_OE				= 1'b0;				// enable ADB output (active LOW)
assign	ADB_SPI_CS			= 1'b1;				// disable serial port interface B

// sinus wave to DA
assign	DA					= o_sine;			// Output sinus wave to DAC A

// Assign 50 kHz Sweep Trigger
assign	sweepTrigger		= GCLKIN;

// Map 50 kHz A-line sweep signal to GPIO[0]
assign	GPIO[0]				= sweepTrigger;

// Receive signal from LabView to record data to DDR2 in GPIO[6]
assign	enableRecording		= GPIO[6];
// Display enable signal from LabView
assign	SEG0_DP				= ~enableRecording;
// Turn off 7-segment displays
assign	SEG0_D				= 1'b0;
assign	SEG1_D				= 1'b0;
assign	SEG1_DP				= 1'b0;
assign 	trigger50kHz		= enableRecording & sweepTrigger;


// Assign 156.25 MHz clock PLL_CLKIN_p to sys_clk
assign	sys_clk				= PLL_CLKIN_p;
assign	FPGA_CLK_A_P		=  sys_clk;
assign	FPGA_CLK_A_N		= ~sys_clk;

//// LED diagnostics
assign	LED[6:4] 			= ~error_data;
//assign	LED[6] 				= ~control_done_read;
assign	LED[3] 				= ~reading_done;
assign	LED[2] 				= ~user_data_available;
//assign	LED[3] 				= ~control_done_write;
assign	LED[1] 				= ~writing_done;
//assign	LED[1] 				= ~user_buffer_full;
assign	LED[0]				= ~error_full;

// Send signal to D6
//assign	GPIO[0]				= user_data_available;
//assign	GPIO[6]				= control_done_read;
//assign	GPIO[1]				= control_go_read;

// Synchronization of sampling with sweep trigger
sample_addressing_custom sample_addressing_custom_inst (
	.clock(ADA_DCO) ,							// input  clock_sig (ADA_DCO)
	.sclr(~trigger50kHz) ,						// input  ~trigger50kHz
	.sample_position(write_RAM_address) ,		// output [10:0] sample_position
	.acq_busy(acq_busy) ,						// output acq_busy
	.acq_done(acq_done) ,						// output acq_done
	.dualMSB_write() ,				// output dualMSB_write
	.dualMSB_read()					// output dualMSB_read
	);

// T flip flop (divides frequency of acq_done by 2)
FlipFlopT	FlipFlopT_inst (
	.clock ( acq_done ),
	.data ( dualMSB_read ),
	.q ( dualMSB_write )
	);

// MSB to read address from internal RAM
assign	dualMSB_read	= ~dualMSB_write;

// 4096 words (16-bit data bus) RAM
RAM	RAM_inst (
	.wraddress ({ dualMSB_write, write_RAM_address }),// Sample position (0-1170)
	.wrclock ( ADA_DCO ),						// Write clock (ADA_DCO or sys_clk????)
	.wren ( acq_busy ),							// acq_busy & ~read_RAM_busy
	.data ( {2'b0, ADA_D} ),					// 16-bit data
	.rdaddress ({ dualMSB_read, read_RAM_address }),// Read adress (read_RAM_address) from NIOS
	.rdclock ( sys_clk ),						// Read clock (sys_clk)
	.q ( RAMdata )								// data read by NIOS
	);

// Ethernet clock PLL
pll_125 pll_125_ins (
	.inclk0(OSC_50_BANK3),
	.c0(enet_refclk_125MHz)
	);

// Generate global reset signal
gen_reset_n	system_gen_reset_n (
	.tx_clk(OSC_50_BANK3),
	.reset_n_in(reset_n),
	.reset_n_out(global_reset_n)
	);

// Generate ethernet reset signal
gen_reset_n	net_gen_reset_n(
	.tx_clk(OSC_50_BANK3),
	.reset_n_in(global_reset_n),
	.reset_n_out(enet_reset_n)
	);
				
// SOPC system with master read and write DDR2 handling
DE4_SOPC DE4_SOPC_inst(
	// 1) global signals:
	.clk_50(OSC_50_BANK3),
	.reset_n(global_reset_n),

`ifndef USE_DDR2_DIMM2
  // the_ddr2
   .aux_scan_clk_from_the_ddr2(),
   .aux_scan_clk_reset_n_from_the_ddr2(),
   .dll_reference_clk_from_the_ddr2(),
   .dqs_delay_ctrl_export_from_the_ddr2(),
   .global_reset_n_to_the_ddr2(reset_n),
   .local_init_done_from_the_ddr2(),
   .local_refresh_ack_from_the_ddr2(),
   .local_wdata_req_from_the_ddr2(),
   .mem_addr_from_the_ddr2(M1_DDR2_addr),
   .mem_ba_from_the_ddr2(M1_DDR2_ba),
   .mem_cas_n_from_the_ddr2(M1_DDR2_cas_n),
   .mem_cke_from_the_ddr2(M1_DDR2_cke),
   .mem_clk_n_to_and_from_the_ddr2(M1_DDR2_clk_n),
   .mem_clk_to_and_from_the_ddr2(M1_DDR2_clk),
   .mem_cs_n_from_the_ddr2(M1_DDR2_cs_n),
   .mem_dm_from_the_ddr2(M1_DDR2_dm),
   .mem_dq_to_and_from_the_ddr2(M1_DDR2_dq),
   .mem_dqs_to_and_from_the_ddr2(M1_DDR2_dqs),
   .mem_dqsn_to_and_from_the_ddr2(M1_DDR2_dqsn),
   .mem_odt_from_the_ddr2(M1_DDR2_odt),
   .mem_ras_n_from_the_ddr2(M1_DDR2_ras_n),
   .mem_we_n_from_the_ddr2(M1_DDR2_we_n),
   .oct_ctl_rs_value_to_the_ddr2(),
   .oct_ctl_rt_value_to_the_ddr2(),
   .reset_phy_clk_n_from_the_ddr2(),
   
  // ddr2 psd i2c
  // NOT NECESSARY WHEN TESING DDR2, ONLY FOR EEPROM
   .out_port_from_the_ddr2_i2c_scl(), 			//M1_DDR2_SCL
   .out_port_from_the_ddr2_i2c_sa(), 			//M1_DDR2_SA
   .bidir_port_to_and_from_the_ddr2_i2c_sda(), 	//M1_DDR2_SDA
   
`else              
	// the_ddr2
	.aux_scan_clk_from_the_ddr2(),
	.aux_scan_clk_reset_n_from_the_ddr2(),
	.dll_reference_clk_from_the_ddr2(),
	.dqs_delay_ctrl_export_from_the_ddr2(),
	.global_reset_n_to_the_ddr2(reset_n),
	.local_init_done_from_the_ddr2(),
	.local_refresh_ack_from_the_ddr2(),
	.local_wdata_req_from_the_ddr2(),
	.mem_addr_from_the_ddr2(M2_DDR2_addr),
	.mem_ba_from_the_ddr2(M2_DDR2_ba),
	.mem_cas_n_from_the_ddr2(M2_DDR2_cas_n),
	.mem_cke_from_the_ddr2(M2_DDR2_cke),
	.mem_clk_n_to_and_from_the_ddr2(M2_DDR2_clk_n),
	.mem_clk_to_and_from_the_ddr2(M2_DDR2_clk),
	.mem_cs_n_from_the_ddr2(M2_DDR2_cs_n),
	.mem_dm_from_the_ddr2(M2_DDR2_dm),
	.mem_dq_to_and_from_the_ddr2(M2_DDR2_dq),
	.mem_dqs_to_and_from_the_ddr2(M2_DDR2_dqs),
	.mem_dqsn_to_and_from_the_ddr2(M2_DDR2_dqsn),
	.mem_odt_from_the_ddr2(M2_DDR2_odt),
	.mem_ras_n_from_the_ddr2(M2_DDR2_ras_n),
	.mem_we_n_from_the_ddr2(M2_DDR2_we_n),
	.oct_ctl_rs_value_to_the_ddr2(),
	.oct_ctl_rt_value_to_the_ddr2(),
	.reset_phy_clk_n_from_the_ddr2(),

	// ddr2 psd i2c
	// NOT NECESSARY WHEN TESING DDR2, ONLY FOR EEPROM
	.out_port_from_the_ddr2_i2c_scl(), 			//M2_DDR2_SCL
	.out_port_from_the_ddr2_i2c_sa(), 			//M2_DDR2_SA
	.bidir_port_to_and_from_the_ddr2_i2c_sda(), //M2_DDR2_SDA       
`endif                   
	
	// clock out
	.ddr2_phy_clk_out (ddr2_phy_clk_out),
	
	// Master Read template
	.control_done_from_the_master_read(control_done_read) ,					// output  
	.control_early_done_from_the_master_read() ,							// output  
	.control_fixed_location_to_the_master_read(0) ,							// input  
	.control_go_to_the_master_read(control_go_read) ,						// input  
	.control_read_base_to_the_master_read(control_read_base) ,				// input [29:0] 
	.control_read_length_to_the_master_read(control_read_length) ,			// input [29:0] 
	.user_buffer_output_data_from_the_master_read(user_buffer_data_read) ,	// output [31:0] 
	.user_data_available_from_the_master_read(user_data_available) ,		// output  
	.user_read_buffer_to_the_master_read(user_read_buffer) ,				// input  
	
	// Master Write template
	.control_done_from_the_master_write(control_done_write) ,				// output  
	.control_fixed_location_to_the_master_write(0) ,						// input  
	.control_go_to_the_master_write(control_go_write) ,						// input  
	.control_write_base_to_the_master_write(control_write_base) ,			// input [29:0] 
	.control_write_length_to_the_master_write(control_write_length) ,		// input [29:0] 
	.user_buffer_full_from_the_master_write(user_buffer_full) ,				// output  
	.user_buffer_input_data_to_the_master_write({224'b0, user_buffer_data_write}) ,	// input [31:0] 
	.user_write_buffer_to_the_master_write(user_write_buffer) 				// input  
	);

// Yields a reset signal 20 ms after cpu reset
//PowerOn_RST PowerOn_RST_inst
//(
//	.clk(OSC_50_BANK3) ,						// input  clk_sig
//	.RSTnCPU(global_reset_n) ,					// input  RSTnCPU_sig
//	.RSTn(reset_power_on) 						// output  RSTn_sig
//);

TestRead TestRead_inst (
	.RSTn(global_reset_n) ,										// input  reset_power_on
	.CLK48MHZ(OSC_50_BANK3) ,									// input  
	.control_go(control_go_read) ,								// output  
	.control_read_base(control_read_base) ,						// output [29:0] 
	.control_read_length(control_read_length) ,					// output [29:0] 
	.control_done(control_done_read) ,							// input  
	.user_buffer_data(user_buffer_data_read[31:0]) ,			// input [31:0] 
	.user_read_buffer(user_read_buffer) ,						// output  
	.user_data_available(user_data_available) ,					// input  
	.addressLastCompleteWrite(address_last_complete_write) ,	// input [29:0] 
	.addressLastCompleteRead(address_last_complete_read) ,		// output [29:0] 
	.readingDone(reading_done) ,								// output  
	.debugOut() ,												// output [31:0] 
	.errorData(error_data) 										// output [2:0] 
	);

TestWrite TestWrite_inst (
	.RSTn(global_reset_n) ,										// input  reset_power_on
	.CLK48MHZ(OSC_50_BANK3) ,									// input  
	.control_go(control_go_write) ,								// output  
	.control_write_base(control_write_base) ,					// output [29:0] 
	.control_write_length(control_write_length) ,				// output [29:0] 
	.control_done(control_done_write) ,							// input  
	.user_buffer_data(user_buffer_data_write) ,					// output [31:0] 
	.user_buffer_full(user_buffer_full) ,						// input  
	.user_write_buffer(user_write_buffer) ,						// output  
	.addressLastCompleteWrite(address_last_complete_write) ,	// output [29:0] 
	.addressLastCompleteRead(address_last_complete_read) ,		// input [29:0] 
	.writingDone(writing_done) ,								// output  
	.debugOut() ,												// output [31:0] 
	.errorFull(error_full) 										// output  
	);

//==============================================================================
// Optional modules
//==============================================================================

// Fan Control
FAN_PWM FAN_PWM_inst (
	.clk(OSC_50_BANK3) ,						// input  OSC_50_BANK3
	.PWM_input(4'hC) ,							// input [3:0] PWM = 4'hC
	.clk_div_out(clk_div_out_sig) ,				// output [7:0] clk_div_out_sig
	.FAN(FAN_CTRL) 								// output FAN_CTRL
	);

// Heartbeat with glowing LED
LED_glow LED_glow_inst (
	.clk(ADA_DCO) ,								// input  clk_div_out_sig[1]
	.LED(LED[7]) 								// output LED_sig
	);

// Generate sinus wave in DAC B to test acquisition
sin400k_st sin400k_st_inst (
	.clk(sys_clk) ,								// input  sys_clk 156.25 MHz clock
	.reset_n(global_reset_n) ,					// input  global_reset_n
	.clken(1'b1) ,								// input  1'b1
	.phi_inc_i(32'd27487791) ,					// input [anglePrec-1:0] @156.25 MHz -> 
												// d10995116 for 400 kHz sinus,
												// d27487791 for 1 MHz.
	.fsin_o(raw_sine) ,							// output [magnitudePrec-1:0] raw_sine
	.out_valid() 								// output  N.C.
	);

// Synchronize DAC A output (sinus wave) with system clock
always @(negedge global_reset_n or posedge sys_clk)
begin
	if (!global_reset_n) begin
		o_sine		<= 14'd0;
	end
	else begin
		// Invert sign bit (MSB) to have offset binary
		o_sine		<= {~raw_sine[13],raw_sine[12:0]};
	end
end

endmodule
