module A_line_acq(
	);
//=======================================================
//  PARAMETER declarations
//=======================================================
parameter

//=======================================================
//  PORT declarations
//=======================================================
input
input
output	reg
//=======================================================
//  REG/WIRE declarations
//=======================================================
reg
wire
//=======================================================
//  Structural coding
//=======================================================	

endmodule