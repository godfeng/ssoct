//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2009 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ad_buf_s1_arbitrator (
                              // inputs:
                               ad_buf_s1_readdata,
                               ad_buf_s1_waitrequest,
                               clk,
                               reset_n,
                               std_2s60_burst_17_downstream_address_to_slave,
                               std_2s60_burst_17_downstream_arbitrationshare,
                               std_2s60_burst_17_downstream_burstcount,
                               std_2s60_burst_17_downstream_latency_counter,
                               std_2s60_burst_17_downstream_read,
                               std_2s60_burst_17_downstream_write,
                               std_2s60_burst_18_downstream_address_to_slave,
                               std_2s60_burst_18_downstream_arbitrationshare,
                               std_2s60_burst_18_downstream_burstcount,
                               std_2s60_burst_18_downstream_latency_counter,
                               std_2s60_burst_18_downstream_read,
                               std_2s60_burst_18_downstream_write,

                              // outputs:
                               ad_buf_s1_address,
                               ad_buf_s1_chipselect_n,
                               ad_buf_s1_read,
                               ad_buf_s1_readdata_from_sa,
                               ad_buf_s1_reset_n,
                               ad_buf_s1_waitrequest_from_sa,
                               d1_ad_buf_s1_end_xfer,
                               std_2s60_burst_17_downstream_granted_ad_buf_s1,
                               std_2s60_burst_17_downstream_qualified_request_ad_buf_s1,
                               std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1,
                               std_2s60_burst_17_downstream_requests_ad_buf_s1,
                               std_2s60_burst_18_downstream_granted_ad_buf_s1,
                               std_2s60_burst_18_downstream_qualified_request_ad_buf_s1,
                               std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1,
                               std_2s60_burst_18_downstream_requests_ad_buf_s1
                            )
;

  output  [ 11: 0] ad_buf_s1_address;
  output           ad_buf_s1_chipselect_n;
  output           ad_buf_s1_read;
  output  [ 31: 0] ad_buf_s1_readdata_from_sa;
  output           ad_buf_s1_reset_n;
  output           ad_buf_s1_waitrequest_from_sa;
  output           d1_ad_buf_s1_end_xfer;
  output           std_2s60_burst_17_downstream_granted_ad_buf_s1;
  output           std_2s60_burst_17_downstream_qualified_request_ad_buf_s1;
  output           std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1;
  output           std_2s60_burst_17_downstream_requests_ad_buf_s1;
  output           std_2s60_burst_18_downstream_granted_ad_buf_s1;
  output           std_2s60_burst_18_downstream_qualified_request_ad_buf_s1;
  output           std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1;
  output           std_2s60_burst_18_downstream_requests_ad_buf_s1;
  input   [ 31: 0] ad_buf_s1_readdata;
  input            ad_buf_s1_waitrequest;
  input            clk;
  input            reset_n;
  input   [ 13: 0] std_2s60_burst_17_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_17_downstream_arbitrationshare;
  input            std_2s60_burst_17_downstream_burstcount;
  input            std_2s60_burst_17_downstream_latency_counter;
  input            std_2s60_burst_17_downstream_read;
  input            std_2s60_burst_17_downstream_write;
  input   [ 13: 0] std_2s60_burst_18_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_18_downstream_arbitrationshare;
  input            std_2s60_burst_18_downstream_burstcount;
  input            std_2s60_burst_18_downstream_latency_counter;
  input            std_2s60_burst_18_downstream_read;
  input            std_2s60_burst_18_downstream_write;

  wire    [ 11: 0] ad_buf_s1_address;
  wire             ad_buf_s1_allgrants;
  wire             ad_buf_s1_allow_new_arb_cycle;
  wire             ad_buf_s1_any_bursting_master_saved_grant;
  wire             ad_buf_s1_any_continuerequest;
  reg     [  1: 0] ad_buf_s1_arb_addend;
  wire             ad_buf_s1_arb_counter_enable;
  reg     [  3: 0] ad_buf_s1_arb_share_counter;
  wire    [  3: 0] ad_buf_s1_arb_share_counter_next_value;
  wire    [  3: 0] ad_buf_s1_arb_share_set_values;
  wire    [  1: 0] ad_buf_s1_arb_winner;
  wire             ad_buf_s1_arbitration_holdoff_internal;
  wire             ad_buf_s1_beginbursttransfer_internal;
  wire             ad_buf_s1_begins_xfer;
  wire             ad_buf_s1_chipselect_n;
  wire    [  3: 0] ad_buf_s1_chosen_master_double_vector;
  wire    [  1: 0] ad_buf_s1_chosen_master_rot_left;
  wire             ad_buf_s1_end_xfer;
  wire             ad_buf_s1_firsttransfer;
  wire    [  1: 0] ad_buf_s1_grant_vector;
  wire             ad_buf_s1_in_a_read_cycle;
  wire             ad_buf_s1_in_a_write_cycle;
  wire    [  1: 0] ad_buf_s1_master_qreq_vector;
  wire             ad_buf_s1_non_bursting_master_requests;
  wire             ad_buf_s1_read;
  wire    [ 31: 0] ad_buf_s1_readdata_from_sa;
  reg              ad_buf_s1_reg_firsttransfer;
  wire             ad_buf_s1_reset_n;
  reg     [  1: 0] ad_buf_s1_saved_chosen_master_vector;
  reg              ad_buf_s1_slavearbiterlockenable;
  wire             ad_buf_s1_slavearbiterlockenable2;
  wire             ad_buf_s1_unreg_firsttransfer;
  wire             ad_buf_s1_waitrequest_from_sa;
  wire             ad_buf_s1_waits_for_read;
  wire             ad_buf_s1_waits_for_write;
  reg              d1_ad_buf_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ad_buf_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_std_2s60_burst_17_downstream_granted_slave_ad_buf_s1;
  reg              last_cycle_std_2s60_burst_18_downstream_granted_slave_ad_buf_s1;
  wire             p1_std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register;
  wire             p1_std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register;
  wire    [ 13: 0] shifted_address_to_ad_buf_s1_from_std_2s60_burst_17_downstream;
  wire    [ 13: 0] shifted_address_to_ad_buf_s1_from_std_2s60_burst_18_downstream;
  wire             std_2s60_burst_17_downstream_arbiterlock;
  wire             std_2s60_burst_17_downstream_arbiterlock2;
  wire             std_2s60_burst_17_downstream_continuerequest;
  wire             std_2s60_burst_17_downstream_granted_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_qualified_request_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1;
  reg              std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register;
  wire             std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register_in;
  wire             std_2s60_burst_17_downstream_requests_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_saved_grant_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_arbiterlock;
  wire             std_2s60_burst_18_downstream_arbiterlock2;
  wire             std_2s60_burst_18_downstream_continuerequest;
  wire             std_2s60_burst_18_downstream_granted_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_qualified_request_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1;
  reg              std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register;
  wire             std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register_in;
  wire             std_2s60_burst_18_downstream_requests_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_saved_grant_ad_buf_s1;
  wire             wait_for_ad_buf_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~ad_buf_s1_end_xfer;
    end


  assign ad_buf_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 | std_2s60_burst_18_downstream_qualified_request_ad_buf_s1));
  //assign ad_buf_s1_readdata_from_sa = ad_buf_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ad_buf_s1_readdata_from_sa = ad_buf_s1_readdata;

  assign std_2s60_burst_17_downstream_requests_ad_buf_s1 = ((1) & (std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write)) & std_2s60_burst_17_downstream_read;
  //assign ad_buf_s1_waitrequest_from_sa = ad_buf_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ad_buf_s1_waitrequest_from_sa = ad_buf_s1_waitrequest;

  //ad_buf_s1_arb_share_counter set values, which is an e_mux
  assign ad_buf_s1_arb_share_set_values = (std_2s60_burst_17_downstream_granted_ad_buf_s1)? std_2s60_burst_17_downstream_arbitrationshare :
    (std_2s60_burst_18_downstream_granted_ad_buf_s1)? std_2s60_burst_18_downstream_arbitrationshare :
    (std_2s60_burst_17_downstream_granted_ad_buf_s1)? std_2s60_burst_17_downstream_arbitrationshare :
    (std_2s60_burst_18_downstream_granted_ad_buf_s1)? std_2s60_burst_18_downstream_arbitrationshare :
    1;

  //ad_buf_s1_non_bursting_master_requests mux, which is an e_mux
  assign ad_buf_s1_non_bursting_master_requests = 0;

  //ad_buf_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ad_buf_s1_any_bursting_master_saved_grant = std_2s60_burst_17_downstream_saved_grant_ad_buf_s1 |
    std_2s60_burst_18_downstream_saved_grant_ad_buf_s1 |
    std_2s60_burst_17_downstream_saved_grant_ad_buf_s1 |
    std_2s60_burst_18_downstream_saved_grant_ad_buf_s1;

  //ad_buf_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ad_buf_s1_arb_share_counter_next_value = ad_buf_s1_firsttransfer ? (ad_buf_s1_arb_share_set_values - 1) : |ad_buf_s1_arb_share_counter ? (ad_buf_s1_arb_share_counter - 1) : 0;

  //ad_buf_s1_allgrants all slave grants, which is an e_mux
  assign ad_buf_s1_allgrants = |ad_buf_s1_grant_vector |
    |ad_buf_s1_grant_vector |
    |ad_buf_s1_grant_vector |
    |ad_buf_s1_grant_vector;

  //ad_buf_s1_end_xfer assignment, which is an e_assign
  assign ad_buf_s1_end_xfer = ~(ad_buf_s1_waits_for_read | ad_buf_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ad_buf_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ad_buf_s1 = ad_buf_s1_end_xfer & (~ad_buf_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ad_buf_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ad_buf_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ad_buf_s1 & ad_buf_s1_allgrants) | (end_xfer_arb_share_counter_term_ad_buf_s1 & ~ad_buf_s1_non_bursting_master_requests);

  //ad_buf_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ad_buf_s1_arb_share_counter <= 0;
      else if (ad_buf_s1_arb_counter_enable)
          ad_buf_s1_arb_share_counter <= ad_buf_s1_arb_share_counter_next_value;
    end


  //ad_buf_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ad_buf_s1_slavearbiterlockenable <= 0;
      else if ((|ad_buf_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ad_buf_s1) | (end_xfer_arb_share_counter_term_ad_buf_s1 & ~ad_buf_s1_non_bursting_master_requests))
          ad_buf_s1_slavearbiterlockenable <= |ad_buf_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_17/downstream ad_buf/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_17_downstream_arbiterlock = ad_buf_s1_slavearbiterlockenable & std_2s60_burst_17_downstream_continuerequest;

  //ad_buf_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ad_buf_s1_slavearbiterlockenable2 = |ad_buf_s1_arb_share_counter_next_value;

  //std_2s60_burst_17/downstream ad_buf/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_17_downstream_arbiterlock2 = ad_buf_s1_slavearbiterlockenable2 & std_2s60_burst_17_downstream_continuerequest;

  //std_2s60_burst_18/downstream ad_buf/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_18_downstream_arbiterlock = ad_buf_s1_slavearbiterlockenable & std_2s60_burst_18_downstream_continuerequest;

  //std_2s60_burst_18/downstream ad_buf/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_18_downstream_arbiterlock2 = ad_buf_s1_slavearbiterlockenable2 & std_2s60_burst_18_downstream_continuerequest;

  //std_2s60_burst_18/downstream granted ad_buf/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_18_downstream_granted_slave_ad_buf_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_18_downstream_granted_slave_ad_buf_s1 <= std_2s60_burst_18_downstream_saved_grant_ad_buf_s1 ? 1 : (ad_buf_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_18_downstream_granted_slave_ad_buf_s1;
    end


  //std_2s60_burst_18_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_18_downstream_continuerequest = last_cycle_std_2s60_burst_18_downstream_granted_slave_ad_buf_s1 & 1;

  //ad_buf_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ad_buf_s1_any_continuerequest = std_2s60_burst_18_downstream_continuerequest |
    std_2s60_burst_17_downstream_continuerequest;

  assign std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 = std_2s60_burst_17_downstream_requests_ad_buf_s1 & ~(std_2s60_burst_18_downstream_arbiterlock);
  //std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register_in = std_2s60_burst_17_downstream_granted_ad_buf_s1 & std_2s60_burst_17_downstream_read & ~ad_buf_s1_waits_for_read;

  //shift register p1 std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register = {std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register, std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register_in};

  //std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register <= p1_std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1, which is an e_mux
  assign std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1 = std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1_shift_register;

  assign std_2s60_burst_18_downstream_requests_ad_buf_s1 = ((1) & (std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write)) & std_2s60_burst_18_downstream_read;
  //std_2s60_burst_17/downstream granted ad_buf/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_17_downstream_granted_slave_ad_buf_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_17_downstream_granted_slave_ad_buf_s1 <= std_2s60_burst_17_downstream_saved_grant_ad_buf_s1 ? 1 : (ad_buf_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_17_downstream_granted_slave_ad_buf_s1;
    end


  //std_2s60_burst_17_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_17_downstream_continuerequest = last_cycle_std_2s60_burst_17_downstream_granted_slave_ad_buf_s1 & 1;

  assign std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 = std_2s60_burst_18_downstream_requests_ad_buf_s1 & ~(std_2s60_burst_17_downstream_arbiterlock);
  //std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register_in = std_2s60_burst_18_downstream_granted_ad_buf_s1 & std_2s60_burst_18_downstream_read & ~ad_buf_s1_waits_for_read;

  //shift register p1 std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register = {std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register, std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register_in};

  //std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register <= p1_std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1, which is an e_mux
  assign std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1 = std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1_shift_register;

  //allow new arb cycle for ad_buf/s1, which is an e_assign
  assign ad_buf_s1_allow_new_arb_cycle = ~std_2s60_burst_17_downstream_arbiterlock & ~std_2s60_burst_18_downstream_arbiterlock;

  //std_2s60_burst_18/downstream assignment into master qualified-requests vector for ad_buf/s1, which is an e_assign
  assign ad_buf_s1_master_qreq_vector[0] = std_2s60_burst_18_downstream_qualified_request_ad_buf_s1;

  //std_2s60_burst_18/downstream grant ad_buf/s1, which is an e_assign
  assign std_2s60_burst_18_downstream_granted_ad_buf_s1 = ad_buf_s1_grant_vector[0];

  //std_2s60_burst_18/downstream saved-grant ad_buf/s1, which is an e_assign
  assign std_2s60_burst_18_downstream_saved_grant_ad_buf_s1 = ad_buf_s1_arb_winner[0];

  //std_2s60_burst_17/downstream assignment into master qualified-requests vector for ad_buf/s1, which is an e_assign
  assign ad_buf_s1_master_qreq_vector[1] = std_2s60_burst_17_downstream_qualified_request_ad_buf_s1;

  //std_2s60_burst_17/downstream grant ad_buf/s1, which is an e_assign
  assign std_2s60_burst_17_downstream_granted_ad_buf_s1 = ad_buf_s1_grant_vector[1];

  //std_2s60_burst_17/downstream saved-grant ad_buf/s1, which is an e_assign
  assign std_2s60_burst_17_downstream_saved_grant_ad_buf_s1 = ad_buf_s1_arb_winner[1];

  //ad_buf/s1 chosen-master double-vector, which is an e_assign
  assign ad_buf_s1_chosen_master_double_vector = {ad_buf_s1_master_qreq_vector, ad_buf_s1_master_qreq_vector} & ({~ad_buf_s1_master_qreq_vector, ~ad_buf_s1_master_qreq_vector} + ad_buf_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign ad_buf_s1_arb_winner = (ad_buf_s1_allow_new_arb_cycle & | ad_buf_s1_grant_vector) ? ad_buf_s1_grant_vector : ad_buf_s1_saved_chosen_master_vector;

  //saved ad_buf_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ad_buf_s1_saved_chosen_master_vector <= 0;
      else if (ad_buf_s1_allow_new_arb_cycle)
          ad_buf_s1_saved_chosen_master_vector <= |ad_buf_s1_grant_vector ? ad_buf_s1_grant_vector : ad_buf_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ad_buf_s1_grant_vector = {(ad_buf_s1_chosen_master_double_vector[1] | ad_buf_s1_chosen_master_double_vector[3]),
    (ad_buf_s1_chosen_master_double_vector[0] | ad_buf_s1_chosen_master_double_vector[2])};

  //ad_buf/s1 chosen master rotated left, which is an e_assign
  assign ad_buf_s1_chosen_master_rot_left = (ad_buf_s1_arb_winner << 1) ? (ad_buf_s1_arb_winner << 1) : 1;

  //ad_buf/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ad_buf_s1_arb_addend <= 1;
      else if (|ad_buf_s1_grant_vector)
          ad_buf_s1_arb_addend <= ad_buf_s1_end_xfer? ad_buf_s1_chosen_master_rot_left : ad_buf_s1_grant_vector;
    end


  //ad_buf_s1_reset_n assignment, which is an e_assign
  assign ad_buf_s1_reset_n = reset_n;

  assign ad_buf_s1_chipselect_n = ~(std_2s60_burst_17_downstream_granted_ad_buf_s1 | std_2s60_burst_18_downstream_granted_ad_buf_s1);
  //ad_buf_s1_firsttransfer first transaction, which is an e_assign
  assign ad_buf_s1_firsttransfer = ad_buf_s1_begins_xfer ? ad_buf_s1_unreg_firsttransfer : ad_buf_s1_reg_firsttransfer;

  //ad_buf_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ad_buf_s1_unreg_firsttransfer = ~(ad_buf_s1_slavearbiterlockenable & ad_buf_s1_any_continuerequest);

  //ad_buf_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ad_buf_s1_reg_firsttransfer <= 1'b1;
      else if (ad_buf_s1_begins_xfer)
          ad_buf_s1_reg_firsttransfer <= ad_buf_s1_unreg_firsttransfer;
    end


  //ad_buf_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ad_buf_s1_beginbursttransfer_internal = ad_buf_s1_begins_xfer;

  //ad_buf_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ad_buf_s1_arbitration_holdoff_internal = ad_buf_s1_begins_xfer & ad_buf_s1_firsttransfer;

  //ad_buf_s1_read assignment, which is an e_mux
  assign ad_buf_s1_read = (std_2s60_burst_17_downstream_granted_ad_buf_s1 & std_2s60_burst_17_downstream_read) | (std_2s60_burst_18_downstream_granted_ad_buf_s1 & std_2s60_burst_18_downstream_read);

  assign shifted_address_to_ad_buf_s1_from_std_2s60_burst_17_downstream = std_2s60_burst_17_downstream_address_to_slave;
  //ad_buf_s1_address mux, which is an e_mux
  assign ad_buf_s1_address = (std_2s60_burst_17_downstream_granted_ad_buf_s1)? (shifted_address_to_ad_buf_s1_from_std_2s60_burst_17_downstream >> 2) :
    (shifted_address_to_ad_buf_s1_from_std_2s60_burst_18_downstream >> 2);

  assign shifted_address_to_ad_buf_s1_from_std_2s60_burst_18_downstream = std_2s60_burst_18_downstream_address_to_slave;
  //d1_ad_buf_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ad_buf_s1_end_xfer <= 1;
      else if (1)
          d1_ad_buf_s1_end_xfer <= ad_buf_s1_end_xfer;
    end


  //ad_buf_s1_waits_for_read in a cycle, which is an e_mux
  assign ad_buf_s1_waits_for_read = ad_buf_s1_in_a_read_cycle & ad_buf_s1_waitrequest_from_sa;

  //ad_buf_s1_in_a_read_cycle assignment, which is an e_assign
  assign ad_buf_s1_in_a_read_cycle = (std_2s60_burst_17_downstream_granted_ad_buf_s1 & std_2s60_burst_17_downstream_read) | (std_2s60_burst_18_downstream_granted_ad_buf_s1 & std_2s60_burst_18_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ad_buf_s1_in_a_read_cycle;

  //ad_buf_s1_waits_for_write in a cycle, which is an e_mux
  assign ad_buf_s1_waits_for_write = ad_buf_s1_in_a_write_cycle & ad_buf_s1_waitrequest_from_sa;

  //ad_buf_s1_in_a_write_cycle assignment, which is an e_assign
  assign ad_buf_s1_in_a_write_cycle = (std_2s60_burst_17_downstream_granted_ad_buf_s1 & std_2s60_burst_17_downstream_write) | (std_2s60_burst_18_downstream_granted_ad_buf_s1 & std_2s60_burst_18_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ad_buf_s1_in_a_write_cycle;

  assign wait_for_ad_buf_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ad_buf/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_17/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_17_downstream_requests_ad_buf_s1 && (std_2s60_burst_17_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_17/downstream drove 0 on its 'arbitrationshare' port while accessing slave ad_buf/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_17/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_17_downstream_requests_ad_buf_s1 && (std_2s60_burst_17_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_17/downstream drove 0 on its 'burstcount' port while accessing slave ad_buf/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_18/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_18_downstream_requests_ad_buf_s1 && (std_2s60_burst_18_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_18/downstream drove 0 on its 'arbitrationshare' port while accessing slave ad_buf/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_18/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_18_downstream_requests_ad_buf_s1 && (std_2s60_burst_18_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_18/downstream drove 0 on its 'burstcount' port while accessing slave ad_buf/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_17_downstream_granted_ad_buf_s1 + std_2s60_burst_18_downstream_granted_ad_buf_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_17_downstream_saved_grant_ad_buf_s1 + std_2s60_burst_18_downstream_saved_grant_ad_buf_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           reset_n,
                                           std_2s60_burst_0_downstream_address_to_slave,
                                           std_2s60_burst_0_downstream_arbitrationshare,
                                           std_2s60_burst_0_downstream_burstcount,
                                           std_2s60_burst_0_downstream_byteenable,
                                           std_2s60_burst_0_downstream_debugaccess,
                                           std_2s60_burst_0_downstream_latency_counter,
                                           std_2s60_burst_0_downstream_read,
                                           std_2s60_burst_0_downstream_write,
                                           std_2s60_burst_0_downstream_writedata,
                                           std_2s60_burst_1_downstream_address_to_slave,
                                           std_2s60_burst_1_downstream_arbitrationshare,
                                           std_2s60_burst_1_downstream_burstcount,
                                           std_2s60_burst_1_downstream_byteenable,
                                           std_2s60_burst_1_downstream_debugaccess,
                                           std_2s60_burst_1_downstream_latency_counter,
                                           std_2s60_burst_1_downstream_read,
                                           std_2s60_burst_1_downstream_write,
                                           std_2s60_burst_1_downstream_writedata,

                                          // outputs:
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer,
                                           std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module,
                                           std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module,
                                           std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module,
                                           std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module,
                                           std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module,
                                           std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module,
                                           std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module,
                                           std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module
                                        )
;

  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  output           std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module;
  output           std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  output           std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;
  output           std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module;
  output           std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;
  output           std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  output           std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;
  output           std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input            reset_n;
  input   [ 10: 0] std_2s60_burst_0_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_0_downstream_arbitrationshare;
  input            std_2s60_burst_0_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_0_downstream_byteenable;
  input            std_2s60_burst_0_downstream_debugaccess;
  input            std_2s60_burst_0_downstream_latency_counter;
  input            std_2s60_burst_0_downstream_read;
  input            std_2s60_burst_0_downstream_write;
  input   [ 31: 0] std_2s60_burst_0_downstream_writedata;
  input   [ 10: 0] std_2s60_burst_1_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_1_downstream_arbitrationshare;
  input            std_2s60_burst_1_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_1_downstream_byteenable;
  input            std_2s60_burst_1_downstream_debugaccess;
  input            std_2s60_burst_1_downstream_latency_counter;
  input            std_2s60_burst_1_downstream_read;
  input            std_2s60_burst_1_downstream_write;
  input   [ 31: 0] std_2s60_burst_1_downstream_writedata;

  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_jtag_debug_module_arb_addend;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg     [  3: 0] cpu_jtag_debug_module_arb_share_counter;
  wire    [  3: 0] cpu_jtag_debug_module_arb_share_counter_next_value;
  wire    [  3: 0] cpu_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_jtag_debug_module_arb_winner;
  wire             cpu_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_std_2s60_burst_0_downstream_granted_slave_cpu_jtag_debug_module;
  reg              last_cycle_std_2s60_burst_1_downstream_granted_slave_cpu_jtag_debug_module;
  wire    [ 10: 0] shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_0_downstream;
  wire    [ 10: 0] shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_1_downstream;
  wire             std_2s60_burst_0_downstream_arbiterlock;
  wire             std_2s60_burst_0_downstream_arbiterlock2;
  wire             std_2s60_burst_0_downstream_continuerequest;
  wire             std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_arbiterlock;
  wire             std_2s60_burst_1_downstream_arbiterlock2;
  wire             std_2s60_burst_1_downstream_continuerequest;
  wire             std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module | std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module = (1) & (std_2s60_burst_0_downstream_read | std_2s60_burst_0_downstream_write);
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_0_downstream_arbitrationshare :
    (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_1_downstream_arbitrationshare :
    (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_0_downstream_arbitrationshare :
    (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_1_downstream_arbitrationshare :
    1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = 0;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module |
    std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module |
    std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module |
    std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = |cpu_jtag_debug_module_grant_vector |
    |cpu_jtag_debug_module_grant_vector |
    |cpu_jtag_debug_module_grant_vector |
    |cpu_jtag_debug_module_grant_vector;

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //std_2s60_burst_0/downstream cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign std_2s60_burst_0_downstream_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & std_2s60_burst_0_downstream_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //std_2s60_burst_0/downstream cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign std_2s60_burst_0_downstream_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & std_2s60_burst_0_downstream_continuerequest;

  //std_2s60_burst_1/downstream cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign std_2s60_burst_1_downstream_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & std_2s60_burst_1_downstream_continuerequest;

  //std_2s60_burst_1/downstream cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign std_2s60_burst_1_downstream_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & std_2s60_burst_1_downstream_continuerequest;

  //std_2s60_burst_1/downstream granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_1_downstream_granted_slave_cpu_jtag_debug_module <= 0;
      else if (1)
          last_cycle_std_2s60_burst_1_downstream_granted_slave_cpu_jtag_debug_module <= std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_1_downstream_granted_slave_cpu_jtag_debug_module;
    end


  //std_2s60_burst_1_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_1_downstream_continuerequest = last_cycle_std_2s60_burst_1_downstream_granted_slave_cpu_jtag_debug_module & 1;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_jtag_debug_module_any_continuerequest = std_2s60_burst_1_downstream_continuerequest |
    std_2s60_burst_0_downstream_continuerequest;

  assign std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module = std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module & ~((std_2s60_burst_0_downstream_read & ((std_2s60_burst_0_downstream_latency_counter != 0))) | std_2s60_burst_1_downstream_arbiterlock);
  //local readdatavalid std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module = std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_0_downstream_read & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_0_downstream_writedata :
    std_2s60_burst_1_downstream_writedata;

  assign std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module = (1) & (std_2s60_burst_1_downstream_read | std_2s60_burst_1_downstream_write);
  //std_2s60_burst_0/downstream granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_0_downstream_granted_slave_cpu_jtag_debug_module <= 0;
      else if (1)
          last_cycle_std_2s60_burst_0_downstream_granted_slave_cpu_jtag_debug_module <= std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_0_downstream_granted_slave_cpu_jtag_debug_module;
    end


  //std_2s60_burst_0_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_0_downstream_continuerequest = last_cycle_std_2s60_burst_0_downstream_granted_slave_cpu_jtag_debug_module & 1;

  assign std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module = std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module & ~((std_2s60_burst_1_downstream_read & ((std_2s60_burst_1_downstream_latency_counter != 0))) | std_2s60_burst_0_downstream_arbiterlock);
  //local readdatavalid std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module = std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_1_downstream_read & ~cpu_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = ~std_2s60_burst_0_downstream_arbiterlock & ~std_2s60_burst_1_downstream_arbiterlock;

  //std_2s60_burst_1/downstream assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[0] = std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module;

  //std_2s60_burst_1/downstream grant cpu/jtag_debug_module, which is an e_assign
  assign std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[0];

  //std_2s60_burst_1/downstream saved-grant cpu/jtag_debug_module, which is an e_assign
  assign std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[0];

  //std_2s60_burst_0/downstream assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[1] = std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module;

  //std_2s60_burst_0/downstream grant cpu/jtag_debug_module, which is an e_assign
  assign std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[1];

  //std_2s60_burst_0/downstream saved-grant cpu/jtag_debug_module, which is an e_assign
  assign std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[1];

  //cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_double_vector = {cpu_jtag_debug_module_master_qreq_vector, cpu_jtag_debug_module_master_qreq_vector} & ({~cpu_jtag_debug_module_master_qreq_vector, ~cpu_jtag_debug_module_master_qreq_vector} + cpu_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_jtag_debug_module_arb_winner = (cpu_jtag_debug_module_allow_new_arb_cycle & | cpu_jtag_debug_module_grant_vector) ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_jtag_debug_module_allow_new_arb_cycle)
          cpu_jtag_debug_module_saved_chosen_master_vector <= |cpu_jtag_debug_module_grant_vector ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_jtag_debug_module_grant_vector = {(cpu_jtag_debug_module_chosen_master_double_vector[1] | cpu_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_jtag_debug_module_chosen_master_double_vector[0] | cpu_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_rot_left = (cpu_jtag_debug_module_arb_winner << 1) ? (cpu_jtag_debug_module_arb_winner << 1) : 1;

  //cpu/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_jtag_debug_module_grant_vector)
          cpu_jtag_debug_module_arb_addend <= cpu_jtag_debug_module_end_xfer? cpu_jtag_debug_module_chosen_master_rot_left : cpu_jtag_debug_module_grant_vector;
    end


  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //assign lhs ~cpu_jtag_debug_module_reset of type reset_n to cpu_jtag_debug_module_reset_n, which is an e_assign
  assign cpu_jtag_debug_module_reset = ~cpu_jtag_debug_module_reset_n;

  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module | std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_jtag_debug_module_arbitration_holdoff_internal = cpu_jtag_debug_module_begins_xfer & cpu_jtag_debug_module_firsttransfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_0_downstream_write) | (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_1_downstream_write);

  assign shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_0_downstream = std_2s60_burst_0_downstream_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? (shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_0_downstream >> 2) :
    (shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_1_downstream >> 2);

  assign shifted_address_to_cpu_jtag_debug_module_from_std_2s60_burst_1_downstream = std_2s60_burst_1_downstream_address_to_slave;
  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else if (1)
          d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_0_downstream_read) | (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_1_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_0_downstream_write) | (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module & std_2s60_burst_1_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_0_downstream_byteenable :
    (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_1_downstream_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_0_downstream_debugaccess :
    (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module)? std_2s60_burst_1_downstream_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module && (std_2s60_burst_0_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end


  //std_2s60_burst_0/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module && (std_2s60_burst_0_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end


  //std_2s60_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module && (std_2s60_burst_1_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end


  //std_2s60_burst_1/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module && (std_2s60_burst_1_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module + std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_0_downstream_saved_grant_cpu_jtag_debug_module + std_2s60_burst_1_downstream_saved_grant_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_burstcount,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_byteenable_std_2s60_burst_3_upstream,
                                     cpu_data_master_granted_std_2s60_burst_10_upstream,
                                     cpu_data_master_granted_std_2s60_burst_11_upstream,
                                     cpu_data_master_granted_std_2s60_burst_12_upstream,
                                     cpu_data_master_granted_std_2s60_burst_13_upstream,
                                     cpu_data_master_granted_std_2s60_burst_14_upstream,
                                     cpu_data_master_granted_std_2s60_burst_16_upstream,
                                     cpu_data_master_granted_std_2s60_burst_17_upstream,
                                     cpu_data_master_granted_std_2s60_burst_1_upstream,
                                     cpu_data_master_granted_std_2s60_burst_3_upstream,
                                     cpu_data_master_granted_std_2s60_burst_5_upstream,
                                     cpu_data_master_granted_std_2s60_burst_7_upstream,
                                     cpu_data_master_granted_std_2s60_burst_9_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_10_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_11_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_12_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_13_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_14_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_16_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_17_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_1_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_3_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_5_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_7_upstream,
                                     cpu_data_master_qualified_request_std_2s60_burst_9_upstream,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_std_2s60_burst_10_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_11_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_12_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_13_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_14_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_16_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_17_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_1_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_3_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_5_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_7_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                     cpu_data_master_read_data_valid_std_2s60_burst_9_upstream,
                                     cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                     cpu_data_master_requests_std_2s60_burst_10_upstream,
                                     cpu_data_master_requests_std_2s60_burst_11_upstream,
                                     cpu_data_master_requests_std_2s60_burst_12_upstream,
                                     cpu_data_master_requests_std_2s60_burst_13_upstream,
                                     cpu_data_master_requests_std_2s60_burst_14_upstream,
                                     cpu_data_master_requests_std_2s60_burst_16_upstream,
                                     cpu_data_master_requests_std_2s60_burst_17_upstream,
                                     cpu_data_master_requests_std_2s60_burst_1_upstream,
                                     cpu_data_master_requests_std_2s60_burst_3_upstream,
                                     cpu_data_master_requests_std_2s60_burst_5_upstream,
                                     cpu_data_master_requests_std_2s60_burst_7_upstream,
                                     cpu_data_master_requests_std_2s60_burst_9_upstream,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     d1_irq_from_the_lan91c111,
                                     d1_std_2s60_burst_10_upstream_end_xfer,
                                     d1_std_2s60_burst_11_upstream_end_xfer,
                                     d1_std_2s60_burst_12_upstream_end_xfer,
                                     d1_std_2s60_burst_13_upstream_end_xfer,
                                     d1_std_2s60_burst_14_upstream_end_xfer,
                                     d1_std_2s60_burst_16_upstream_end_xfer,
                                     d1_std_2s60_burst_17_upstream_end_xfer,
                                     d1_std_2s60_burst_1_upstream_end_xfer,
                                     d1_std_2s60_burst_3_upstream_end_xfer,
                                     d1_std_2s60_burst_5_upstream_end_xfer,
                                     d1_std_2s60_burst_7_upstream_end_xfer,
                                     d1_std_2s60_burst_9_upstream_end_xfer,
                                     high_res_timer_s1_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     reset_n,
                                     std_2s60_burst_10_upstream_readdata_from_sa,
                                     std_2s60_burst_10_upstream_waitrequest_from_sa,
                                     std_2s60_burst_11_upstream_readdata_from_sa,
                                     std_2s60_burst_11_upstream_waitrequest_from_sa,
                                     std_2s60_burst_12_upstream_readdata_from_sa,
                                     std_2s60_burst_12_upstream_waitrequest_from_sa,
                                     std_2s60_burst_13_upstream_readdata_from_sa,
                                     std_2s60_burst_13_upstream_waitrequest_from_sa,
                                     std_2s60_burst_14_upstream_readdata_from_sa,
                                     std_2s60_burst_14_upstream_waitrequest_from_sa,
                                     std_2s60_burst_16_upstream_readdata_from_sa,
                                     std_2s60_burst_16_upstream_waitrequest_from_sa,
                                     std_2s60_burst_17_upstream_readdata_from_sa,
                                     std_2s60_burst_17_upstream_waitrequest_from_sa,
                                     std_2s60_burst_1_upstream_readdata_from_sa,
                                     std_2s60_burst_1_upstream_waitrequest_from_sa,
                                     std_2s60_burst_3_upstream_readdata_from_sa,
                                     std_2s60_burst_3_upstream_waitrequest_from_sa,
                                     std_2s60_burst_5_upstream_readdata_from_sa,
                                     std_2s60_burst_5_upstream_waitrequest_from_sa,
                                     std_2s60_burst_7_upstream_readdata_from_sa,
                                     std_2s60_burst_7_upstream_waitrequest_from_sa,
                                     std_2s60_burst_9_upstream_readdata_from_sa,
                                     std_2s60_burst_9_upstream_waitrequest_from_sa,
                                     sys_clk_timer_s1_irq_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_dbs_address,
                                     cpu_data_master_dbs_write_8,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 25: 0] cpu_data_master_address_to_slave;
  output  [  1: 0] cpu_data_master_dbs_address;
  output  [  7: 0] cpu_data_master_dbs_write_8;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input            clk;
  input   [ 25: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_byteenable_std_2s60_burst_3_upstream;
  input            cpu_data_master_granted_std_2s60_burst_10_upstream;
  input            cpu_data_master_granted_std_2s60_burst_11_upstream;
  input            cpu_data_master_granted_std_2s60_burst_12_upstream;
  input            cpu_data_master_granted_std_2s60_burst_13_upstream;
  input            cpu_data_master_granted_std_2s60_burst_14_upstream;
  input            cpu_data_master_granted_std_2s60_burst_16_upstream;
  input            cpu_data_master_granted_std_2s60_burst_17_upstream;
  input            cpu_data_master_granted_std_2s60_burst_1_upstream;
  input            cpu_data_master_granted_std_2s60_burst_3_upstream;
  input            cpu_data_master_granted_std_2s60_burst_5_upstream;
  input            cpu_data_master_granted_std_2s60_burst_7_upstream;
  input            cpu_data_master_granted_std_2s60_burst_9_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_10_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_11_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_12_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_13_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_14_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_16_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_17_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_1_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_3_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_5_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_7_upstream;
  input            cpu_data_master_qualified_request_std_2s60_burst_9_upstream;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_requests_std_2s60_burst_10_upstream;
  input            cpu_data_master_requests_std_2s60_burst_11_upstream;
  input            cpu_data_master_requests_std_2s60_burst_12_upstream;
  input            cpu_data_master_requests_std_2s60_burst_13_upstream;
  input            cpu_data_master_requests_std_2s60_burst_14_upstream;
  input            cpu_data_master_requests_std_2s60_burst_16_upstream;
  input            cpu_data_master_requests_std_2s60_burst_17_upstream;
  input            cpu_data_master_requests_std_2s60_burst_1_upstream;
  input            cpu_data_master_requests_std_2s60_burst_3_upstream;
  input            cpu_data_master_requests_std_2s60_burst_5_upstream;
  input            cpu_data_master_requests_std_2s60_burst_7_upstream;
  input            cpu_data_master_requests_std_2s60_burst_9_upstream;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            d1_irq_from_the_lan91c111;
  input            d1_std_2s60_burst_10_upstream_end_xfer;
  input            d1_std_2s60_burst_11_upstream_end_xfer;
  input            d1_std_2s60_burst_12_upstream_end_xfer;
  input            d1_std_2s60_burst_13_upstream_end_xfer;
  input            d1_std_2s60_burst_14_upstream_end_xfer;
  input            d1_std_2s60_burst_16_upstream_end_xfer;
  input            d1_std_2s60_burst_17_upstream_end_xfer;
  input            d1_std_2s60_burst_1_upstream_end_xfer;
  input            d1_std_2s60_burst_3_upstream_end_xfer;
  input            d1_std_2s60_burst_5_upstream_end_xfer;
  input            d1_std_2s60_burst_7_upstream_end_xfer;
  input            d1_std_2s60_burst_9_upstream_end_xfer;
  input            high_res_timer_s1_irq_from_sa;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_10_upstream_readdata_from_sa;
  input            std_2s60_burst_10_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_11_upstream_readdata_from_sa;
  input            std_2s60_burst_11_upstream_waitrequest_from_sa;
  input   [ 15: 0] std_2s60_burst_12_upstream_readdata_from_sa;
  input            std_2s60_burst_12_upstream_waitrequest_from_sa;
  input   [  7: 0] std_2s60_burst_13_upstream_readdata_from_sa;
  input            std_2s60_burst_13_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_14_upstream_readdata_from_sa;
  input            std_2s60_burst_14_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_16_upstream_readdata_from_sa;
  input            std_2s60_burst_16_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_17_upstream_readdata_from_sa;
  input            std_2s60_burst_17_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_1_upstream_readdata_from_sa;
  input            std_2s60_burst_1_upstream_waitrequest_from_sa;
  input   [  7: 0] std_2s60_burst_3_upstream_readdata_from_sa;
  input            std_2s60_burst_3_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_5_upstream_readdata_from_sa;
  input            std_2s60_burst_5_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_7_upstream_readdata_from_sa;
  input            std_2s60_burst_7_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_9_upstream_readdata_from_sa;
  input            std_2s60_burst_9_upstream_waitrequest_from_sa;
  input            sys_clk_timer_s1_irq_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 25: 0] cpu_data_master_address_last_time;
  wire    [ 25: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_burstcount_last_time;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_data_master_dbs_address;
  wire    [  1: 0] cpu_data_master_dbs_increment;
  reg     [  1: 0] cpu_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_data_master_dbs_rdv_counter_inc;
  wire    [  7: 0] cpu_data_master_dbs_write_8;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg              cpu_data_master_latency_counter;
  wire    [  1: 0] cpu_data_master_next_dbs_rdv_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [  7: 0] dbs_latent_8_reg_segment_0;
  reg     [  7: 0] dbs_latent_8_reg_segment_1;
  reg     [  7: 0] dbs_latent_8_reg_segment_2;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_data_master_latency_counter;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_2;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_std_2s60_burst_1_upstream | ~cpu_data_master_requests_std_2s60_burst_1_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_1_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_1_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_1_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_1_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_10_upstream | ~cpu_data_master_requests_std_2s60_burst_10_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_10_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_10_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_10_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_10_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_11_upstream | ~cpu_data_master_requests_std_2s60_burst_11_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_11_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_11_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_11_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_11_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_12_upstream | ~cpu_data_master_requests_std_2s60_burst_12_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_12_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_12_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_12_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_12_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_13_upstream | ~cpu_data_master_requests_std_2s60_burst_13_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_13_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_13_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_13_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_13_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_data_master_qualified_request_std_2s60_burst_14_upstream | ~cpu_data_master_requests_std_2s60_burst_14_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_14_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_14_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_14_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_14_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_16_upstream | ~cpu_data_master_requests_std_2s60_burst_16_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_16_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_16_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_16_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_16_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_17_upstream | ~cpu_data_master_requests_std_2s60_burst_17_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_17_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_17_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_17_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_17_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_3_upstream | ~cpu_data_master_requests_std_2s60_burst_3_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_3_upstream | ~cpu_data_master_read | (1 & ~std_2s60_burst_3_upstream_waitrequest_from_sa & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_std_2s60_burst_3_upstream | ~cpu_data_master_write | (1 & ~std_2s60_burst_3_upstream_waitrequest_from_sa & (cpu_data_master_dbs_address[1] & cpu_data_master_dbs_address[0]) & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_5_upstream | ~cpu_data_master_requests_std_2s60_burst_5_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_5_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_5_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_5_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_5_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_data_master_qualified_request_std_2s60_burst_7_upstream | ~cpu_data_master_requests_std_2s60_burst_7_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_7_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_7_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_7_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_7_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_std_2s60_burst_9_upstream | ~cpu_data_master_requests_std_2s60_burst_9_upstream) & ((~cpu_data_master_qualified_request_std_2s60_burst_9_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_9_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_std_2s60_burst_9_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~std_2s60_burst_9_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    high_res_timer_s1_irq_from_sa,
    d1_irq_from_the_lan91c111,
    jtag_uart_avalon_jtag_slave_irq_from_sa,
    sys_clk_timer_s1_irq_from_sa};

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[25 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else if (1)
          cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_std_2s60_burst_1_upstream |
    cpu_data_master_granted_std_2s60_burst_10_upstream |
    cpu_data_master_granted_std_2s60_burst_11_upstream |
    cpu_data_master_granted_std_2s60_burst_12_upstream |
    cpu_data_master_granted_std_2s60_burst_13_upstream |
    cpu_data_master_granted_std_2s60_burst_14_upstream |
    cpu_data_master_granted_std_2s60_burst_16_upstream |
    cpu_data_master_granted_std_2s60_burst_17_upstream |
    cpu_data_master_granted_std_2s60_burst_3_upstream |
    cpu_data_master_granted_std_2s60_burst_5_upstream |
    cpu_data_master_granted_std_2s60_burst_7_upstream |
    cpu_data_master_granted_std_2s60_burst_9_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_std_2s60_burst_1_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_10_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_11_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_12_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_13_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_14_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_16_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_17_upstream |
    (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream & dbs_rdv_counter_overflow) |
    cpu_data_master_read_data_valid_std_2s60_burst_5_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_7_upstream |
    cpu_data_master_read_data_valid_std_2s60_burst_9_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_1_upstream}} | std_2s60_burst_1_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_10_upstream}} | std_2s60_burst_10_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_11_upstream}} | std_2s60_burst_11_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_12_upstream}} | std_2s60_burst_12_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_13_upstream}} | std_2s60_burst_13_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_14_upstream}} | std_2s60_burst_14_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_16_upstream}} | std_2s60_burst_16_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_17_upstream}} | std_2s60_burst_17_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_3_upstream}} | {std_2s60_burst_3_upstream_readdata_from_sa[7 : 0],
    dbs_latent_8_reg_segment_2,
    dbs_latent_8_reg_segment_1,
    dbs_latent_8_reg_segment_0}) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_5_upstream}} | std_2s60_burst_5_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_7_upstream}} | std_2s60_burst_7_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_std_2s60_burst_9_upstream}} | std_2s60_burst_9_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else if (1)
          cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //input to latent dbs-8 stored 0, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_0 = std_2s60_burst_3_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_data_master_dbs_rdv_counter[1 : 0]) == 0))
          dbs_latent_8_reg_segment_0 <= p1_dbs_latent_8_reg_segment_0;
    end


  //input to latent dbs-8 stored 1, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_1 = std_2s60_burst_3_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_1 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_data_master_dbs_rdv_counter[1 : 0]) == 1))
          dbs_latent_8_reg_segment_1 <= p1_dbs_latent_8_reg_segment_1;
    end


  //input to latent dbs-8 stored 2, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_2 = std_2s60_burst_3_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_2 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_data_master_dbs_rdv_counter[1 : 0]) == 2))
          dbs_latent_8_reg_segment_2 <= p1_dbs_latent_8_reg_segment_2;
    end


  //mux write dbs 2, which is an e_mux
  assign cpu_data_master_dbs_write_8 = ((cpu_data_master_dbs_address[1 : 0] == 0))? cpu_data_master_writedata[7 : 0] :
    ((cpu_data_master_dbs_address[1 : 0] == 1))? cpu_data_master_writedata[15 : 8] :
    ((cpu_data_master_dbs_address[1 : 0] == 2))? cpu_data_master_writedata[23 : 16] :
    cpu_data_master_writedata[31 : 24];

  //dbs count increment, which is an e_mux
  assign cpu_data_master_dbs_increment = (cpu_data_master_requests_std_2s60_burst_3_upstream)? 1 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_data_master_dbs_address + cpu_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_data_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_data_master_next_dbs_rdv_counter = cpu_data_master_dbs_rdv_counter + cpu_data_master_dbs_rdv_counter_inc;

  //cpu_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_data_master_dbs_rdv_counter_inc = 1;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_data_master_read_data_valid_std_2s60_burst_3_upstream;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_data_master_dbs_rdv_counter <= cpu_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_data_master_dbs_rdv_counter[1] & ~cpu_data_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_read & 0 & 1 & ~std_2s60_burst_3_upstream_waitrequest_from_sa) |
    (cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_write & 1 & 1 & ~std_2s60_burst_3_upstream_waitrequest_from_sa);


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else if (1)
          cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_burstcount_last_time <= 0;
      else if (1)
          cpu_data_master_burstcount_last_time <= cpu_data_master_burstcount;
    end


  //cpu_data_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_burstcount != cpu_data_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_data_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else if (1)
          cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else if (1)
          cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else if (1)
          cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else if (1)
          cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_burstcount,
                                            cpu_instruction_master_granted_std_2s60_burst_0_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_15_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_18_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_2_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_4_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_6_upstream,
                                            cpu_instruction_master_granted_std_2s60_burst_8_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream,
                                            cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream,
                                            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                            cpu_instruction_master_requests_std_2s60_burst_0_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_15_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_18_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_2_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_4_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_6_upstream,
                                            cpu_instruction_master_requests_std_2s60_burst_8_upstream,
                                            d1_std_2s60_burst_0_upstream_end_xfer,
                                            d1_std_2s60_burst_15_upstream_end_xfer,
                                            d1_std_2s60_burst_18_upstream_end_xfer,
                                            d1_std_2s60_burst_2_upstream_end_xfer,
                                            d1_std_2s60_burst_4_upstream_end_xfer,
                                            d1_std_2s60_burst_6_upstream_end_xfer,
                                            d1_std_2s60_burst_8_upstream_end_xfer,
                                            reset_n,
                                            std_2s60_burst_0_upstream_readdata_from_sa,
                                            std_2s60_burst_0_upstream_waitrequest_from_sa,
                                            std_2s60_burst_15_upstream_readdata_from_sa,
                                            std_2s60_burst_15_upstream_waitrequest_from_sa,
                                            std_2s60_burst_18_upstream_readdata_from_sa,
                                            std_2s60_burst_18_upstream_waitrequest_from_sa,
                                            std_2s60_burst_2_upstream_readdata_from_sa,
                                            std_2s60_burst_2_upstream_waitrequest_from_sa,
                                            std_2s60_burst_4_upstream_readdata_from_sa,
                                            std_2s60_burst_4_upstream_waitrequest_from_sa,
                                            std_2s60_burst_6_upstream_readdata_from_sa,
                                            std_2s60_burst_6_upstream_waitrequest_from_sa,
                                            std_2s60_burst_8_upstream_readdata_from_sa,
                                            std_2s60_burst_8_upstream_waitrequest_from_sa,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_dbs_address,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 25: 0] cpu_instruction_master_address_to_slave;
  output  [  1: 0] cpu_instruction_master_dbs_address;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_granted_std_2s60_burst_0_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_15_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_18_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_2_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_4_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_6_upstream;
  input            cpu_instruction_master_granted_std_2s60_burst_8_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream;
  input            cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            cpu_instruction_master_requests_std_2s60_burst_0_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_15_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_18_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_2_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_4_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_6_upstream;
  input            cpu_instruction_master_requests_std_2s60_burst_8_upstream;
  input            d1_std_2s60_burst_0_upstream_end_xfer;
  input            d1_std_2s60_burst_15_upstream_end_xfer;
  input            d1_std_2s60_burst_18_upstream_end_xfer;
  input            d1_std_2s60_burst_2_upstream_end_xfer;
  input            d1_std_2s60_burst_4_upstream_end_xfer;
  input            d1_std_2s60_burst_6_upstream_end_xfer;
  input            d1_std_2s60_burst_8_upstream_end_xfer;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_0_upstream_readdata_from_sa;
  input            std_2s60_burst_0_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_15_upstream_readdata_from_sa;
  input            std_2s60_burst_15_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_18_upstream_readdata_from_sa;
  input            std_2s60_burst_18_upstream_waitrequest_from_sa;
  input   [  7: 0] std_2s60_burst_2_upstream_readdata_from_sa;
  input            std_2s60_burst_2_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_4_upstream_readdata_from_sa;
  input            std_2s60_burst_4_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_6_upstream_readdata_from_sa;
  input            std_2s60_burst_6_upstream_waitrequest_from_sa;
  input   [ 31: 0] std_2s60_burst_8_upstream_readdata_from_sa;
  input            std_2s60_burst_8_upstream_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 25: 0] cpu_instruction_master_address_last_time;
  wire    [ 25: 0] cpu_instruction_master_address_to_slave;
  reg     [  3: 0] cpu_instruction_master_burstcount_last_time;
  reg     [  1: 0] cpu_instruction_master_dbs_address;
  wire    [  1: 0] cpu_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  wire    [  1: 0] cpu_instruction_master_next_dbs_rdv_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [  7: 0] dbs_latent_8_reg_segment_0;
  reg     [  7: 0] dbs_latent_8_reg_segment_1;
  reg     [  7: 0] dbs_latent_8_reg_segment_2;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_instruction_master_latency_counter;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_latent_8_reg_segment_2;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream | ~cpu_instruction_master_requests_std_2s60_burst_0_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_0_upstream_waitrequest_from_sa & (cpu_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream | ~cpu_instruction_master_requests_std_2s60_burst_15_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_15_upstream_waitrequest_from_sa & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream | ~cpu_instruction_master_requests_std_2s60_burst_18_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_18_upstream_waitrequest_from_sa & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream | ~cpu_instruction_master_requests_std_2s60_burst_2_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream | ~cpu_instruction_master_read | (1 & ~std_2s60_burst_2_upstream_waitrequest_from_sa & cpu_instruction_master_read))) & 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream | ~cpu_instruction_master_requests_std_2s60_burst_4_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_4_upstream_waitrequest_from_sa & (cpu_instruction_master_read))));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream | ~cpu_instruction_master_requests_std_2s60_burst_6_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_6_upstream_waitrequest_from_sa & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream | ~cpu_instruction_master_requests_std_2s60_burst_8_upstream) & ((~cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream | ~(cpu_instruction_master_read) | (1 & ~std_2s60_burst_8_upstream_waitrequest_from_sa & (cpu_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = cpu_instruction_master_address[25 : 0];

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else if (1)
          cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_std_2s60_burst_0_upstream |
    cpu_instruction_master_granted_std_2s60_burst_15_upstream |
    cpu_instruction_master_granted_std_2s60_burst_18_upstream |
    cpu_instruction_master_granted_std_2s60_burst_2_upstream |
    cpu_instruction_master_granted_std_2s60_burst_4_upstream |
    cpu_instruction_master_granted_std_2s60_burst_6_upstream |
    cpu_instruction_master_granted_std_2s60_burst_8_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream |
    cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream |
    cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream |
    (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream & dbs_rdv_counter_overflow) |
    cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream |
    cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream |
    cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream}} | std_2s60_burst_0_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream}} | std_2s60_burst_15_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream}} | std_2s60_burst_18_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream}} | {std_2s60_burst_2_upstream_readdata_from_sa[7 : 0],
    dbs_latent_8_reg_segment_2,
    dbs_latent_8_reg_segment_1,
    dbs_latent_8_reg_segment_0}) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream}} | std_2s60_burst_4_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream}} | std_2s60_burst_6_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream}} | std_2s60_burst_8_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else if (1)
          cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //input to latent dbs-8 stored 0, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_0 = std_2s60_burst_2_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_instruction_master_dbs_rdv_counter[1 : 0]) == 0))
          dbs_latent_8_reg_segment_0 <= p1_dbs_latent_8_reg_segment_0;
    end


  //input to latent dbs-8 stored 1, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_1 = std_2s60_burst_2_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_1 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_instruction_master_dbs_rdv_counter[1 : 0]) == 1))
          dbs_latent_8_reg_segment_1 <= p1_dbs_latent_8_reg_segment_1;
    end


  //input to latent dbs-8 stored 2, which is an e_mux
  assign p1_dbs_latent_8_reg_segment_2 = std_2s60_burst_2_upstream_readdata_from_sa;

  //dbs register for latent dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_8_reg_segment_2 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_instruction_master_dbs_rdv_counter[1 : 0]) == 2))
          dbs_latent_8_reg_segment_2 <= p1_dbs_latent_8_reg_segment_2;
    end


  //dbs count increment, which is an e_mux
  assign cpu_instruction_master_dbs_increment = (cpu_instruction_master_requests_std_2s60_burst_2_upstream)? 1 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_instruction_master_dbs_address + cpu_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_instruction_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_instruction_master_next_dbs_rdv_counter = cpu_instruction_master_dbs_rdv_counter + cpu_instruction_master_dbs_rdv_counter_inc;

  //cpu_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_instruction_master_dbs_rdv_counter_inc = 1;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_instruction_master_dbs_rdv_counter <= cpu_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_instruction_master_dbs_rdv_counter[1] & ~cpu_instruction_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = cpu_instruction_master_granted_std_2s60_burst_2_upstream & cpu_instruction_master_read & 0 & 1 & ~std_2s60_burst_2_upstream_waitrequest_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else if (1)
          cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_burstcount_last_time <= 0;
      else if (1)
          cpu_instruction_master_burstcount_last_time <= cpu_instruction_master_burstcount;
    end


  //cpu_instruction_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_burstcount != cpu_instruction_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else if (1)
          cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_bus_avalon_slave_arbitrator (
                                               // inputs:
                                                clk,
                                                reset_n,
                                                std_2s60_burst_2_downstream_address_to_slave,
                                                std_2s60_burst_2_downstream_arbitrationshare,
                                                std_2s60_burst_2_downstream_burstcount,
                                                std_2s60_burst_2_downstream_byteenable,
                                                std_2s60_burst_2_downstream_latency_counter,
                                                std_2s60_burst_2_downstream_read,
                                                std_2s60_burst_2_downstream_write,
                                                std_2s60_burst_2_downstream_writedata,
                                                std_2s60_burst_3_downstream_address_to_slave,
                                                std_2s60_burst_3_downstream_arbitrationshare,
                                                std_2s60_burst_3_downstream_burstcount,
                                                std_2s60_burst_3_downstream_byteenable,
                                                std_2s60_burst_3_downstream_latency_counter,
                                                std_2s60_burst_3_downstream_read,
                                                std_2s60_burst_3_downstream_write,
                                                std_2s60_burst_3_downstream_writedata,

                                               // outputs:
                                                d1_ext_flash_bus_avalon_slave_end_xfer,
                                                ext_flash_bus_address,
                                                ext_flash_bus_data,
                                                ext_flash_bus_readn,
                                                ext_flash_s1_wait_counter_eq_0,
                                                incoming_ext_flash_bus_data_with_Xs_converted_to_0,
                                                select_n_to_the_ext_flash,
                                                std_2s60_burst_2_downstream_granted_ext_flash_s1,
                                                std_2s60_burst_2_downstream_qualified_request_ext_flash_s1,
                                                std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1,
                                                std_2s60_burst_2_downstream_requests_ext_flash_s1,
                                                std_2s60_burst_3_downstream_granted_ext_flash_s1,
                                                std_2s60_burst_3_downstream_qualified_request_ext_flash_s1,
                                                std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1,
                                                std_2s60_burst_3_downstream_requests_ext_flash_s1,
                                                write_n_to_the_ext_flash
                                             )
;

  output           d1_ext_flash_bus_avalon_slave_end_xfer;
  output  [ 23: 0] ext_flash_bus_address;
  inout   [  7: 0] ext_flash_bus_data;
  output           ext_flash_bus_readn;
  output           ext_flash_s1_wait_counter_eq_0;
  output  [  7: 0] incoming_ext_flash_bus_data_with_Xs_converted_to_0;
  output           select_n_to_the_ext_flash;
  output           std_2s60_burst_2_downstream_granted_ext_flash_s1;
  output           std_2s60_burst_2_downstream_qualified_request_ext_flash_s1;
  output           std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1;
  output           std_2s60_burst_2_downstream_requests_ext_flash_s1;
  output           std_2s60_burst_3_downstream_granted_ext_flash_s1;
  output           std_2s60_burst_3_downstream_qualified_request_ext_flash_s1;
  output           std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1;
  output           std_2s60_burst_3_downstream_requests_ext_flash_s1;
  output           write_n_to_the_ext_flash;
  input            clk;
  input            reset_n;
  input   [ 23: 0] std_2s60_burst_2_downstream_address_to_slave;
  input   [  5: 0] std_2s60_burst_2_downstream_arbitrationshare;
  input            std_2s60_burst_2_downstream_burstcount;
  input            std_2s60_burst_2_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_2_downstream_latency_counter;
  input            std_2s60_burst_2_downstream_read;
  input            std_2s60_burst_2_downstream_write;
  input   [  7: 0] std_2s60_burst_2_downstream_writedata;
  input   [ 23: 0] std_2s60_burst_3_downstream_address_to_slave;
  input   [  5: 0] std_2s60_burst_3_downstream_arbitrationshare;
  input            std_2s60_burst_3_downstream_burstcount;
  input            std_2s60_burst_3_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_3_downstream_latency_counter;
  input            std_2s60_burst_3_downstream_read;
  input            std_2s60_burst_3_downstream_write;
  input   [  7: 0] std_2s60_burst_3_downstream_writedata;

  reg              d1_ext_flash_bus_avalon_slave_end_xfer;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [  7: 0] d1_outgoing_ext_flash_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave;
  reg     [ 23: 0] ext_flash_bus_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             ext_flash_bus_avalon_slave_allgrants;
  wire             ext_flash_bus_avalon_slave_allow_new_arb_cycle;
  wire             ext_flash_bus_avalon_slave_any_bursting_master_saved_grant;
  wire             ext_flash_bus_avalon_slave_any_continuerequest;
  reg     [  1: 0] ext_flash_bus_avalon_slave_arb_addend;
  wire             ext_flash_bus_avalon_slave_arb_counter_enable;
  reg     [  5: 0] ext_flash_bus_avalon_slave_arb_share_counter;
  wire    [  5: 0] ext_flash_bus_avalon_slave_arb_share_counter_next_value;
  wire    [  5: 0] ext_flash_bus_avalon_slave_arb_share_set_values;
  wire    [  1: 0] ext_flash_bus_avalon_slave_arb_winner;
  wire             ext_flash_bus_avalon_slave_arbitration_holdoff_internal;
  wire             ext_flash_bus_avalon_slave_beginbursttransfer_internal;
  wire             ext_flash_bus_avalon_slave_begins_xfer;
  wire    [  3: 0] ext_flash_bus_avalon_slave_chosen_master_double_vector;
  wire    [  1: 0] ext_flash_bus_avalon_slave_chosen_master_rot_left;
  wire             ext_flash_bus_avalon_slave_end_xfer;
  wire             ext_flash_bus_avalon_slave_firsttransfer;
  wire    [  1: 0] ext_flash_bus_avalon_slave_grant_vector;
  wire    [  1: 0] ext_flash_bus_avalon_slave_master_qreq_vector;
  wire             ext_flash_bus_avalon_slave_non_bursting_master_requests;
  wire             ext_flash_bus_avalon_slave_read_pending;
  reg              ext_flash_bus_avalon_slave_reg_firsttransfer;
  reg     [  1: 0] ext_flash_bus_avalon_slave_saved_chosen_master_vector;
  reg              ext_flash_bus_avalon_slave_slavearbiterlockenable;
  wire             ext_flash_bus_avalon_slave_slavearbiterlockenable2;
  wire             ext_flash_bus_avalon_slave_unreg_firsttransfer;
  wire             ext_flash_bus_avalon_slave_write_pending;
  wire    [  7: 0] ext_flash_bus_data;
  reg              ext_flash_bus_readn /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire    [  5: 0] ext_flash_s1_counter_load_value;
  wire             ext_flash_s1_in_a_read_cycle;
  wire             ext_flash_s1_in_a_write_cycle;
  wire             ext_flash_s1_pretend_byte_enable;
  reg     [  5: 0] ext_flash_s1_wait_counter;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire             ext_flash_s1_waits_for_read;
  wire             ext_flash_s1_waits_for_write;
  wire             ext_flash_s1_with_write_latency;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [  7: 0] incoming_ext_flash_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_ext_flash_bus_data_bit_0_is_x;
  wire             incoming_ext_flash_bus_data_bit_1_is_x;
  wire             incoming_ext_flash_bus_data_bit_2_is_x;
  wire             incoming_ext_flash_bus_data_bit_3_is_x;
  wire             incoming_ext_flash_bus_data_bit_4_is_x;
  wire             incoming_ext_flash_bus_data_bit_5_is_x;
  wire             incoming_ext_flash_bus_data_bit_6_is_x;
  wire             incoming_ext_flash_bus_data_bit_7_is_x;
  wire    [  7: 0] incoming_ext_flash_bus_data_with_Xs_converted_to_0;
  reg              last_cycle_std_2s60_burst_2_downstream_granted_slave_ext_flash_s1;
  reg              last_cycle_std_2s60_burst_3_downstream_granted_slave_ext_flash_s1;
  wire    [  7: 0] outgoing_ext_flash_bus_data;
  wire    [ 23: 0] p1_ext_flash_bus_address;
  wire             p1_ext_flash_bus_readn;
  wire             p1_select_n_to_the_ext_flash;
  wire    [  1: 0] p1_std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register;
  wire             p1_write_n_to_the_ext_flash;
  reg              select_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             std_2s60_burst_2_downstream_arbiterlock;
  wire             std_2s60_burst_2_downstream_arbiterlock2;
  wire             std_2s60_burst_2_downstream_continuerequest;
  wire             std_2s60_burst_2_downstream_granted_ext_flash_s1;
  wire             std_2s60_burst_2_downstream_qualified_request_ext_flash_s1;
  wire             std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1;
  reg     [  1: 0] std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register;
  wire             std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register_in;
  wire             std_2s60_burst_2_downstream_requests_ext_flash_s1;
  wire             std_2s60_burst_2_downstream_saved_grant_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_arbiterlock;
  wire             std_2s60_burst_3_downstream_arbiterlock2;
  wire             std_2s60_burst_3_downstream_continuerequest;
  wire             std_2s60_burst_3_downstream_granted_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_qualified_request_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1;
  reg     [  1: 0] std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register;
  wire             std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register_in;
  wire             std_2s60_burst_3_downstream_requests_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_saved_grant_ext_flash_s1;
  wire             time_to_write;
  wire             wait_for_ext_flash_s1_counter;
  reg              write_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~ext_flash_bus_avalon_slave_end_xfer;
    end


  assign ext_flash_bus_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 | std_2s60_burst_3_downstream_qualified_request_ext_flash_s1));
  assign std_2s60_burst_2_downstream_requests_ext_flash_s1 = (1) & (std_2s60_burst_2_downstream_read | std_2s60_burst_2_downstream_write);
  //~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_flash <= ~0;
      else if (1)
          select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end


  assign ext_flash_bus_avalon_slave_write_pending = 0;
  //ext_flash_bus/avalon_slave read pending calc, which is an e_assign
  assign ext_flash_bus_avalon_slave_read_pending = 0;

  //ext_flash_bus_avalon_slave_arb_share_counter set values, which is an e_mux
  assign ext_flash_bus_avalon_slave_arb_share_set_values = (std_2s60_burst_2_downstream_granted_ext_flash_s1)? std_2s60_burst_2_downstream_arbitrationshare :
    (std_2s60_burst_3_downstream_granted_ext_flash_s1)? std_2s60_burst_3_downstream_arbitrationshare :
    (std_2s60_burst_2_downstream_granted_ext_flash_s1)? std_2s60_burst_2_downstream_arbitrationshare :
    (std_2s60_burst_3_downstream_granted_ext_flash_s1)? std_2s60_burst_3_downstream_arbitrationshare :
    1;

  //ext_flash_bus_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign ext_flash_bus_avalon_slave_non_bursting_master_requests = 0;

  //ext_flash_bus_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign ext_flash_bus_avalon_slave_any_bursting_master_saved_grant = std_2s60_burst_2_downstream_saved_grant_ext_flash_s1 |
    std_2s60_burst_3_downstream_saved_grant_ext_flash_s1 |
    std_2s60_burst_2_downstream_saved_grant_ext_flash_s1 |
    std_2s60_burst_3_downstream_saved_grant_ext_flash_s1;

  //ext_flash_bus_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign ext_flash_bus_avalon_slave_arb_share_counter_next_value = ext_flash_bus_avalon_slave_firsttransfer ? (ext_flash_bus_avalon_slave_arb_share_set_values - 1) : |ext_flash_bus_avalon_slave_arb_share_counter ? (ext_flash_bus_avalon_slave_arb_share_counter - 1) : 0;

  //ext_flash_bus_avalon_slave_allgrants all slave grants, which is an e_mux
  assign ext_flash_bus_avalon_slave_allgrants = |ext_flash_bus_avalon_slave_grant_vector |
    |ext_flash_bus_avalon_slave_grant_vector |
    |ext_flash_bus_avalon_slave_grant_vector |
    |ext_flash_bus_avalon_slave_grant_vector;

  //ext_flash_bus_avalon_slave_end_xfer assignment, which is an e_assign
  assign ext_flash_bus_avalon_slave_end_xfer = ~(ext_flash_s1_waits_for_read | ext_flash_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave = ext_flash_bus_avalon_slave_end_xfer & (~ext_flash_bus_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ext_flash_bus_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign ext_flash_bus_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave & ext_flash_bus_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave & ~ext_flash_bus_avalon_slave_non_bursting_master_requests);

  //ext_flash_bus_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_avalon_slave_arb_share_counter <= 0;
      else if (ext_flash_bus_avalon_slave_arb_counter_enable)
          ext_flash_bus_avalon_slave_arb_share_counter <= ext_flash_bus_avalon_slave_arb_share_counter_next_value;
    end


  //ext_flash_bus_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|ext_flash_bus_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave) | (end_xfer_arb_share_counter_term_ext_flash_bus_avalon_slave & ~ext_flash_bus_avalon_slave_non_bursting_master_requests))
          ext_flash_bus_avalon_slave_slavearbiterlockenable <= |ext_flash_bus_avalon_slave_arb_share_counter_next_value;
    end


  //std_2s60_burst_2/downstream ext_flash_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_2_downstream_arbiterlock = ext_flash_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_2_downstream_continuerequest;

  //ext_flash_bus_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ext_flash_bus_avalon_slave_slavearbiterlockenable2 = |ext_flash_bus_avalon_slave_arb_share_counter_next_value;

  //std_2s60_burst_2/downstream ext_flash_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_2_downstream_arbiterlock2 = ext_flash_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_2_downstream_continuerequest;

  //std_2s60_burst_3/downstream ext_flash_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_3_downstream_arbiterlock = ext_flash_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_3_downstream_continuerequest;

  //std_2s60_burst_3/downstream ext_flash_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_3_downstream_arbiterlock2 = ext_flash_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_3_downstream_continuerequest;

  //std_2s60_burst_3/downstream granted ext_flash/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_3_downstream_granted_slave_ext_flash_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_3_downstream_granted_slave_ext_flash_s1 <= std_2s60_burst_3_downstream_saved_grant_ext_flash_s1 ? 1 : (ext_flash_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_3_downstream_granted_slave_ext_flash_s1;
    end


  //std_2s60_burst_3_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_3_downstream_continuerequest = last_cycle_std_2s60_burst_3_downstream_granted_slave_ext_flash_s1 & 1;

  //ext_flash_bus_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ext_flash_bus_avalon_slave_any_continuerequest = std_2s60_burst_3_downstream_continuerequest |
    std_2s60_burst_2_downstream_continuerequest;

  assign std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 = std_2s60_burst_2_downstream_requests_ext_flash_s1 & ~((std_2s60_burst_2_downstream_read & (ext_flash_bus_avalon_slave_write_pending | (ext_flash_bus_avalon_slave_read_pending))) | ((ext_flash_bus_avalon_slave_read_pending) & std_2s60_burst_2_downstream_write) | std_2s60_burst_3_downstream_arbiterlock);
  //std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register_in = std_2s60_burst_2_downstream_granted_ext_flash_s1 & std_2s60_burst_2_downstream_read & ~ext_flash_s1_waits_for_read;

  //shift register p1 std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register = {std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register, std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register_in};

  //std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register <= p1_std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1, which is an e_mux
  assign std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1 = std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1_shift_register[1];

  //ext_flash_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_ext_flash_bus_data <= 0;
      else if (1)
          incoming_ext_flash_bus_data <= ext_flash_bus_data;
    end


  //ext_flash_s1_with_write_latency assignment, which is an e_assign
  assign ext_flash_s1_with_write_latency = in_a_write_cycle & (std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 | std_2s60_burst_3_downstream_qualified_request_ext_flash_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (ext_flash_s1_with_write_latency)? 1 :
    (ext_flash_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_ext_flash_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_ext_flash_bus_data <= 0;
      else if (1)
          d1_outgoing_ext_flash_bus_data <= outgoing_ext_flash_bus_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else if (1)
          d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_ext_flash_bus_data tristate driver, which is an e_assign
  assign ext_flash_bus_data = (d1_in_a_write_cycle)? d1_outgoing_ext_flash_bus_data:{8{1'bz}};

  //outgoing_ext_flash_bus_data mux, which is an e_mux
  assign outgoing_ext_flash_bus_data = (std_2s60_burst_2_downstream_granted_ext_flash_s1)? std_2s60_burst_2_downstream_writedata :
    std_2s60_burst_3_downstream_writedata;

  assign std_2s60_burst_3_downstream_requests_ext_flash_s1 = (1) & (std_2s60_burst_3_downstream_read | std_2s60_burst_3_downstream_write);
  //std_2s60_burst_2/downstream granted ext_flash/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_2_downstream_granted_slave_ext_flash_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_2_downstream_granted_slave_ext_flash_s1 <= std_2s60_burst_2_downstream_saved_grant_ext_flash_s1 ? 1 : (ext_flash_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_2_downstream_granted_slave_ext_flash_s1;
    end


  //std_2s60_burst_2_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_2_downstream_continuerequest = last_cycle_std_2s60_burst_2_downstream_granted_slave_ext_flash_s1 & 1;

  assign std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 = std_2s60_burst_3_downstream_requests_ext_flash_s1 & ~((std_2s60_burst_3_downstream_read & (ext_flash_bus_avalon_slave_write_pending | (ext_flash_bus_avalon_slave_read_pending))) | ((ext_flash_bus_avalon_slave_read_pending) & std_2s60_burst_3_downstream_write) | std_2s60_burst_2_downstream_arbiterlock);
  //std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register_in = std_2s60_burst_3_downstream_granted_ext_flash_s1 & std_2s60_burst_3_downstream_read & ~ext_flash_s1_waits_for_read;

  //shift register p1 std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register = {std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register, std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register_in};

  //std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register <= p1_std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1, which is an e_mux
  assign std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1 = std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1_shift_register[1];

  //allow new arb cycle for ext_flash_bus/avalon_slave, which is an e_assign
  assign ext_flash_bus_avalon_slave_allow_new_arb_cycle = ~std_2s60_burst_2_downstream_arbiterlock & ~std_2s60_burst_3_downstream_arbiterlock;

  //std_2s60_burst_3/downstream assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  assign ext_flash_bus_avalon_slave_master_qreq_vector[0] = std_2s60_burst_3_downstream_qualified_request_ext_flash_s1;

  //std_2s60_burst_3/downstream grant ext_flash/s1, which is an e_assign
  assign std_2s60_burst_3_downstream_granted_ext_flash_s1 = ext_flash_bus_avalon_slave_grant_vector[0];

  //std_2s60_burst_3/downstream saved-grant ext_flash/s1, which is an e_assign
  assign std_2s60_burst_3_downstream_saved_grant_ext_flash_s1 = ext_flash_bus_avalon_slave_arb_winner[0];

  //std_2s60_burst_2/downstream assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  assign ext_flash_bus_avalon_slave_master_qreq_vector[1] = std_2s60_burst_2_downstream_qualified_request_ext_flash_s1;

  //std_2s60_burst_2/downstream grant ext_flash/s1, which is an e_assign
  assign std_2s60_burst_2_downstream_granted_ext_flash_s1 = ext_flash_bus_avalon_slave_grant_vector[1];

  //std_2s60_burst_2/downstream saved-grant ext_flash/s1, which is an e_assign
  assign std_2s60_burst_2_downstream_saved_grant_ext_flash_s1 = ext_flash_bus_avalon_slave_arb_winner[1];

  //ext_flash_bus/avalon_slave chosen-master double-vector, which is an e_assign
  assign ext_flash_bus_avalon_slave_chosen_master_double_vector = {ext_flash_bus_avalon_slave_master_qreq_vector, ext_flash_bus_avalon_slave_master_qreq_vector} & ({~ext_flash_bus_avalon_slave_master_qreq_vector, ~ext_flash_bus_avalon_slave_master_qreq_vector} + ext_flash_bus_avalon_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign ext_flash_bus_avalon_slave_arb_winner = (ext_flash_bus_avalon_slave_allow_new_arb_cycle & | ext_flash_bus_avalon_slave_grant_vector) ? ext_flash_bus_avalon_slave_grant_vector : ext_flash_bus_avalon_slave_saved_chosen_master_vector;

  //saved ext_flash_bus_avalon_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_avalon_slave_saved_chosen_master_vector <= 0;
      else if (ext_flash_bus_avalon_slave_allow_new_arb_cycle)
          ext_flash_bus_avalon_slave_saved_chosen_master_vector <= |ext_flash_bus_avalon_slave_grant_vector ? ext_flash_bus_avalon_slave_grant_vector : ext_flash_bus_avalon_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ext_flash_bus_avalon_slave_grant_vector = {(ext_flash_bus_avalon_slave_chosen_master_double_vector[1] | ext_flash_bus_avalon_slave_chosen_master_double_vector[3]),
    (ext_flash_bus_avalon_slave_chosen_master_double_vector[0] | ext_flash_bus_avalon_slave_chosen_master_double_vector[2])};

  //ext_flash_bus/avalon_slave chosen master rotated left, which is an e_assign
  assign ext_flash_bus_avalon_slave_chosen_master_rot_left = (ext_flash_bus_avalon_slave_arb_winner << 1) ? (ext_flash_bus_avalon_slave_arb_winner << 1) : 1;

  //ext_flash_bus/avalon_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_avalon_slave_arb_addend <= 1;
      else if (|ext_flash_bus_avalon_slave_grant_vector)
          ext_flash_bus_avalon_slave_arb_addend <= ext_flash_bus_avalon_slave_end_xfer? ext_flash_bus_avalon_slave_chosen_master_rot_left : ext_flash_bus_avalon_slave_grant_vector;
    end


  assign p1_select_n_to_the_ext_flash = ~(std_2s60_burst_2_downstream_granted_ext_flash_s1 | std_2s60_burst_3_downstream_granted_ext_flash_s1);
  //ext_flash_bus_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign ext_flash_bus_avalon_slave_firsttransfer = ext_flash_bus_avalon_slave_begins_xfer ? ext_flash_bus_avalon_slave_unreg_firsttransfer : ext_flash_bus_avalon_slave_reg_firsttransfer;

  //ext_flash_bus_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign ext_flash_bus_avalon_slave_unreg_firsttransfer = ~(ext_flash_bus_avalon_slave_slavearbiterlockenable & ext_flash_bus_avalon_slave_any_continuerequest);

  //ext_flash_bus_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (ext_flash_bus_avalon_slave_begins_xfer)
          ext_flash_bus_avalon_slave_reg_firsttransfer <= ext_flash_bus_avalon_slave_unreg_firsttransfer;
    end


  //ext_flash_bus_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ext_flash_bus_avalon_slave_beginbursttransfer_internal = ext_flash_bus_avalon_slave_begins_xfer;

  //ext_flash_bus_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ext_flash_bus_avalon_slave_arbitration_holdoff_internal = ext_flash_bus_avalon_slave_begins_xfer & ext_flash_bus_avalon_slave_firsttransfer;

  //~ext_flash_bus_readn of type read to ~p1_ext_flash_bus_readn, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_readn <= ~0;
      else if (1)
          ext_flash_bus_readn <= p1_ext_flash_bus_readn;
    end


  //~p1_ext_flash_bus_readn assignment, which is an e_mux
  assign p1_ext_flash_bus_readn = ~(((std_2s60_burst_2_downstream_granted_ext_flash_s1 & std_2s60_burst_2_downstream_read) | (std_2s60_burst_3_downstream_granted_ext_flash_s1 & std_2s60_burst_3_downstream_read))& ~ext_flash_bus_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter < 26));

  //~write_n_to_the_ext_flash of type write to ~p1_write_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_n_to_the_ext_flash <= ~0;
      else if (1)
          write_n_to_the_ext_flash <= p1_write_n_to_the_ext_flash;
    end


  //~p1_write_n_to_the_ext_flash assignment, which is an e_mux
  assign p1_write_n_to_the_ext_flash = ~(((std_2s60_burst_2_downstream_granted_ext_flash_s1 & std_2s60_burst_2_downstream_write) | (std_2s60_burst_3_downstream_granted_ext_flash_s1 & std_2s60_burst_3_downstream_write)) & ~ext_flash_bus_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter >= 6) & (ext_flash_s1_wait_counter < 32) & ext_flash_s1_pretend_byte_enable);

  //ext_flash_bus_address of type address to p1_ext_flash_bus_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_bus_address <= 0;
      else if (1)
          ext_flash_bus_address <= p1_ext_flash_bus_address;
    end


  //p1_ext_flash_bus_address mux, which is an e_mux
  assign p1_ext_flash_bus_address = (std_2s60_burst_2_downstream_granted_ext_flash_s1)? std_2s60_burst_2_downstream_address_to_slave :
    std_2s60_burst_3_downstream_address_to_slave;

  //d1_ext_flash_bus_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ext_flash_bus_avalon_slave_end_xfer <= 1;
      else if (1)
          d1_ext_flash_bus_avalon_slave_end_xfer <= ext_flash_bus_avalon_slave_end_xfer;
    end


  //ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_read = ext_flash_s1_in_a_read_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_read_cycle = (std_2s60_burst_2_downstream_granted_ext_flash_s1 & std_2s60_burst_2_downstream_read) | (std_2s60_burst_3_downstream_granted_ext_flash_s1 & std_2s60_burst_3_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ext_flash_s1_in_a_read_cycle;

  //ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_write = ext_flash_s1_in_a_write_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_write_cycle = (std_2s60_burst_2_downstream_granted_ext_flash_s1 & std_2s60_burst_2_downstream_write) | (std_2s60_burst_3_downstream_granted_ext_flash_s1 & std_2s60_burst_3_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ext_flash_s1_in_a_write_cycle;

  assign ext_flash_s1_wait_counter_eq_0 = ext_flash_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_s1_wait_counter <= 0;
      else if (1)
          ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end


  assign ext_flash_s1_counter_load_value = ((ext_flash_s1_in_a_read_cycle & ext_flash_bus_avalon_slave_begins_xfer))? 32 :
    ((ext_flash_s1_in_a_write_cycle & ext_flash_bus_avalon_slave_begins_xfer))? 38 :
    (~ext_flash_s1_wait_counter_eq_0)? ext_flash_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_flash_s1_counter = ext_flash_bus_avalon_slave_begins_xfer | ~ext_flash_s1_wait_counter_eq_0;
  //ext_flash_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  assign ext_flash_s1_pretend_byte_enable = (std_2s60_burst_2_downstream_granted_ext_flash_s1)? std_2s60_burst_2_downstream_byteenable :
    (std_2s60_burst_3_downstream_granted_ext_flash_s1)? std_2s60_burst_3_downstream_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //incoming_ext_flash_bus_data_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_0_is_x = ^(incoming_ext_flash_bus_data[0]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[0] = incoming_ext_flash_bus_data_bit_0_is_x ? 1'b0 : incoming_ext_flash_bus_data[0];

  //incoming_ext_flash_bus_data_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_1_is_x = ^(incoming_ext_flash_bus_data[1]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[1] = incoming_ext_flash_bus_data_bit_1_is_x ? 1'b0 : incoming_ext_flash_bus_data[1];

  //incoming_ext_flash_bus_data_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_2_is_x = ^(incoming_ext_flash_bus_data[2]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[2] = incoming_ext_flash_bus_data_bit_2_is_x ? 1'b0 : incoming_ext_flash_bus_data[2];

  //incoming_ext_flash_bus_data_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_3_is_x = ^(incoming_ext_flash_bus_data[3]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[3] = incoming_ext_flash_bus_data_bit_3_is_x ? 1'b0 : incoming_ext_flash_bus_data[3];

  //incoming_ext_flash_bus_data_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_4_is_x = ^(incoming_ext_flash_bus_data[4]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[4] = incoming_ext_flash_bus_data_bit_4_is_x ? 1'b0 : incoming_ext_flash_bus_data[4];

  //incoming_ext_flash_bus_data_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_5_is_x = ^(incoming_ext_flash_bus_data[5]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[5] = incoming_ext_flash_bus_data_bit_5_is_x ? 1'b0 : incoming_ext_flash_bus_data[5];

  //incoming_ext_flash_bus_data_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_6_is_x = ^(incoming_ext_flash_bus_data[6]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[6] = incoming_ext_flash_bus_data_bit_6_is_x ? 1'b0 : incoming_ext_flash_bus_data[6];

  //incoming_ext_flash_bus_data_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_ext_flash_bus_data_bit_7_is_x = ^(incoming_ext_flash_bus_data[7]) === 1'bx;

  //Crush incoming_ext_flash_bus_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0[7] = incoming_ext_flash_bus_data_bit_7_is_x ? 1'b0 : incoming_ext_flash_bus_data[7];

  //ext_flash/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_2_downstream_requests_ext_flash_s1 && (std_2s60_burst_2_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave ext_flash/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_2/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_2_downstream_requests_ext_flash_s1 && (std_2s60_burst_2_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave ext_flash/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_3_downstream_requests_ext_flash_s1 && (std_2s60_burst_3_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave ext_flash/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_3/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_3_downstream_requests_ext_flash_s1 && (std_2s60_burst_3_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave ext_flash/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_2_downstream_granted_ext_flash_s1 + std_2s60_burst_3_downstream_granted_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_2_downstream_saved_grant_ext_flash_s1 + std_2s60_burst_3_downstream_saved_grant_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_ext_flash_bus_data_with_Xs_converted_to_0 = incoming_ext_flash_bus_data;
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_bus_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_bus_avalon_slave_arbitrator (
                                             // inputs:
                                              clk,
                                              irq_from_the_lan91c111,
                                              reset_n,
                                              std_2s60_burst_4_downstream_address_to_slave,
                                              std_2s60_burst_4_downstream_arbitrationshare,
                                              std_2s60_burst_4_downstream_burstcount,
                                              std_2s60_burst_4_downstream_byteenable,
                                              std_2s60_burst_4_downstream_latency_counter,
                                              std_2s60_burst_4_downstream_nativeaddress,
                                              std_2s60_burst_4_downstream_read,
                                              std_2s60_burst_4_downstream_write,
                                              std_2s60_burst_4_downstream_writedata,
                                              std_2s60_burst_5_downstream_address_to_slave,
                                              std_2s60_burst_5_downstream_arbitrationshare,
                                              std_2s60_burst_5_downstream_burstcount,
                                              std_2s60_burst_5_downstream_byteenable,
                                              std_2s60_burst_5_downstream_latency_counter,
                                              std_2s60_burst_5_downstream_nativeaddress,
                                              std_2s60_burst_5_downstream_read,
                                              std_2s60_burst_5_downstream_write,
                                              std_2s60_burst_5_downstream_writedata,
                                              std_2s60_burst_8_downstream_address_to_slave,
                                              std_2s60_burst_8_downstream_arbitrationshare,
                                              std_2s60_burst_8_downstream_burstcount,
                                              std_2s60_burst_8_downstream_byteenable,
                                              std_2s60_burst_8_downstream_latency_counter,
                                              std_2s60_burst_8_downstream_nativeaddress,
                                              std_2s60_burst_8_downstream_read,
                                              std_2s60_burst_8_downstream_write,
                                              std_2s60_burst_8_downstream_writedata,
                                              std_2s60_burst_9_downstream_address_to_slave,
                                              std_2s60_burst_9_downstream_arbitrationshare,
                                              std_2s60_burst_9_downstream_burstcount,
                                              std_2s60_burst_9_downstream_byteenable,
                                              std_2s60_burst_9_downstream_latency_counter,
                                              std_2s60_burst_9_downstream_nativeaddress,
                                              std_2s60_burst_9_downstream_read,
                                              std_2s60_burst_9_downstream_write,
                                              std_2s60_burst_9_downstream_writedata,

                                             // outputs:
                                              be_n_to_the_ext_ram,
                                              d1_ext_ram_bus_avalon_slave_end_xfer,
                                              d1_irq_from_the_lan91c111,
                                              ext_ram_bus_address,
                                              ext_ram_bus_byteenablen,
                                              ext_ram_bus_data,
                                              ext_ram_s1_wait_counter_eq_0,
                                              incoming_ext_ram_bus_data,
                                              ior_n_to_the_lan91c111,
                                              iow_n_to_the_lan91c111,
                                              lan91c111_s1_wait_counter_eq_0,
                                              read_n_to_the_ext_ram,
                                              reset_to_the_lan91c111,
                                              select_n_to_the_ext_ram,
                                              std_2s60_burst_4_downstream_granted_ext_ram_s1,
                                              std_2s60_burst_4_downstream_granted_lan91c111_s1,
                                              std_2s60_burst_4_downstream_qualified_request_ext_ram_s1,
                                              std_2s60_burst_4_downstream_qualified_request_lan91c111_s1,
                                              std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1,
                                              std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1,
                                              std_2s60_burst_4_downstream_requests_ext_ram_s1,
                                              std_2s60_burst_4_downstream_requests_lan91c111_s1,
                                              std_2s60_burst_5_downstream_granted_ext_ram_s1,
                                              std_2s60_burst_5_downstream_granted_lan91c111_s1,
                                              std_2s60_burst_5_downstream_qualified_request_ext_ram_s1,
                                              std_2s60_burst_5_downstream_qualified_request_lan91c111_s1,
                                              std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1,
                                              std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1,
                                              std_2s60_burst_5_downstream_requests_ext_ram_s1,
                                              std_2s60_burst_5_downstream_requests_lan91c111_s1,
                                              std_2s60_burst_8_downstream_granted_ext_ram_s1,
                                              std_2s60_burst_8_downstream_granted_lan91c111_s1,
                                              std_2s60_burst_8_downstream_qualified_request_ext_ram_s1,
                                              std_2s60_burst_8_downstream_qualified_request_lan91c111_s1,
                                              std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1,
                                              std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1,
                                              std_2s60_burst_8_downstream_requests_ext_ram_s1,
                                              std_2s60_burst_8_downstream_requests_lan91c111_s1,
                                              std_2s60_burst_9_downstream_granted_ext_ram_s1,
                                              std_2s60_burst_9_downstream_granted_lan91c111_s1,
                                              std_2s60_burst_9_downstream_qualified_request_ext_ram_s1,
                                              std_2s60_burst_9_downstream_qualified_request_lan91c111_s1,
                                              std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1,
                                              std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1,
                                              std_2s60_burst_9_downstream_requests_ext_ram_s1,
                                              std_2s60_burst_9_downstream_requests_lan91c111_s1,
                                              write_n_to_the_ext_ram
                                           )
;

  output  [  3: 0] be_n_to_the_ext_ram;
  output           d1_ext_ram_bus_avalon_slave_end_xfer;
  output           d1_irq_from_the_lan91c111;
  output  [ 19: 0] ext_ram_bus_address;
  output  [  3: 0] ext_ram_bus_byteenablen;
  inout   [ 31: 0] ext_ram_bus_data;
  output           ext_ram_s1_wait_counter_eq_0;
  output  [ 31: 0] incoming_ext_ram_bus_data;
  output           ior_n_to_the_lan91c111;
  output           iow_n_to_the_lan91c111;
  output           lan91c111_s1_wait_counter_eq_0;
  output           read_n_to_the_ext_ram;
  output           reset_to_the_lan91c111;
  output           select_n_to_the_ext_ram;
  output           std_2s60_burst_4_downstream_granted_ext_ram_s1;
  output           std_2s60_burst_4_downstream_granted_lan91c111_s1;
  output           std_2s60_burst_4_downstream_qualified_request_ext_ram_s1;
  output           std_2s60_burst_4_downstream_qualified_request_lan91c111_s1;
  output           std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1;
  output           std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1;
  output           std_2s60_burst_4_downstream_requests_ext_ram_s1;
  output           std_2s60_burst_4_downstream_requests_lan91c111_s1;
  output           std_2s60_burst_5_downstream_granted_ext_ram_s1;
  output           std_2s60_burst_5_downstream_granted_lan91c111_s1;
  output           std_2s60_burst_5_downstream_qualified_request_ext_ram_s1;
  output           std_2s60_burst_5_downstream_qualified_request_lan91c111_s1;
  output           std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1;
  output           std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1;
  output           std_2s60_burst_5_downstream_requests_ext_ram_s1;
  output           std_2s60_burst_5_downstream_requests_lan91c111_s1;
  output           std_2s60_burst_8_downstream_granted_ext_ram_s1;
  output           std_2s60_burst_8_downstream_granted_lan91c111_s1;
  output           std_2s60_burst_8_downstream_qualified_request_ext_ram_s1;
  output           std_2s60_burst_8_downstream_qualified_request_lan91c111_s1;
  output           std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1;
  output           std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1;
  output           std_2s60_burst_8_downstream_requests_ext_ram_s1;
  output           std_2s60_burst_8_downstream_requests_lan91c111_s1;
  output           std_2s60_burst_9_downstream_granted_ext_ram_s1;
  output           std_2s60_burst_9_downstream_granted_lan91c111_s1;
  output           std_2s60_burst_9_downstream_qualified_request_ext_ram_s1;
  output           std_2s60_burst_9_downstream_qualified_request_lan91c111_s1;
  output           std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1;
  output           std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1;
  output           std_2s60_burst_9_downstream_requests_ext_ram_s1;
  output           std_2s60_burst_9_downstream_requests_lan91c111_s1;
  output           write_n_to_the_ext_ram;
  input            clk;
  input            irq_from_the_lan91c111;
  input            reset_n;
  input   [ 19: 0] std_2s60_burst_4_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_4_downstream_arbitrationshare;
  input            std_2s60_burst_4_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_4_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_4_downstream_latency_counter;
  input   [ 19: 0] std_2s60_burst_4_downstream_nativeaddress;
  input            std_2s60_burst_4_downstream_read;
  input            std_2s60_burst_4_downstream_write;
  input   [ 31: 0] std_2s60_burst_4_downstream_writedata;
  input   [ 19: 0] std_2s60_burst_5_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_5_downstream_arbitrationshare;
  input            std_2s60_burst_5_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_5_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_5_downstream_latency_counter;
  input   [ 19: 0] std_2s60_burst_5_downstream_nativeaddress;
  input            std_2s60_burst_5_downstream_read;
  input            std_2s60_burst_5_downstream_write;
  input   [ 31: 0] std_2s60_burst_5_downstream_writedata;
  input   [ 15: 0] std_2s60_burst_8_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_8_downstream_arbitrationshare;
  input            std_2s60_burst_8_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_8_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_8_downstream_latency_counter;
  input   [ 15: 0] std_2s60_burst_8_downstream_nativeaddress;
  input            std_2s60_burst_8_downstream_read;
  input            std_2s60_burst_8_downstream_write;
  input   [ 31: 0] std_2s60_burst_8_downstream_writedata;
  input   [ 15: 0] std_2s60_burst_9_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_9_downstream_arbitrationshare;
  input            std_2s60_burst_9_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_9_downstream_byteenable;
  input   [  1: 0] std_2s60_burst_9_downstream_latency_counter;
  input   [ 15: 0] std_2s60_burst_9_downstream_nativeaddress;
  input            std_2s60_burst_9_downstream_read;
  input            std_2s60_burst_9_downstream_write;
  input   [ 31: 0] std_2s60_burst_9_downstream_writedata;

  reg     [  3: 0] be_n_to_the_ext_ram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_ext_ram_bus_avalon_slave_end_xfer;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg              d1_irq_from_the_lan91c111;
  reg     [ 31: 0] d1_outgoing_ext_ram_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave;
  reg     [ 19: 0] ext_ram_bus_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             ext_ram_bus_avalon_slave_allgrants;
  wire             ext_ram_bus_avalon_slave_allow_new_arb_cycle;
  wire             ext_ram_bus_avalon_slave_any_bursting_master_saved_grant;
  wire             ext_ram_bus_avalon_slave_any_continuerequest;
  reg     [  7: 0] ext_ram_bus_avalon_slave_arb_addend;
  wire             ext_ram_bus_avalon_slave_arb_counter_enable;
  reg     [  3: 0] ext_ram_bus_avalon_slave_arb_share_counter;
  wire    [  3: 0] ext_ram_bus_avalon_slave_arb_share_counter_next_value;
  wire    [  3: 0] ext_ram_bus_avalon_slave_arb_share_set_values;
  wire    [  7: 0] ext_ram_bus_avalon_slave_arb_winner;
  wire             ext_ram_bus_avalon_slave_arbitration_holdoff_internal;
  wire             ext_ram_bus_avalon_slave_beginbursttransfer_internal;
  wire             ext_ram_bus_avalon_slave_begins_xfer;
  wire    [ 15: 0] ext_ram_bus_avalon_slave_chosen_master_double_vector;
  wire    [  7: 0] ext_ram_bus_avalon_slave_chosen_master_rot_left;
  wire             ext_ram_bus_avalon_slave_end_xfer;
  wire             ext_ram_bus_avalon_slave_firsttransfer;
  wire    [  7: 0] ext_ram_bus_avalon_slave_grant_vector;
  wire    [  7: 0] ext_ram_bus_avalon_slave_master_qreq_vector;
  wire             ext_ram_bus_avalon_slave_non_bursting_master_requests;
  wire             ext_ram_bus_avalon_slave_read_pending;
  reg              ext_ram_bus_avalon_slave_reg_firsttransfer;
  reg     [  7: 0] ext_ram_bus_avalon_slave_saved_chosen_master_vector;
  reg              ext_ram_bus_avalon_slave_slavearbiterlockenable;
  wire             ext_ram_bus_avalon_slave_slavearbiterlockenable2;
  wire             ext_ram_bus_avalon_slave_unreg_firsttransfer;
  wire             ext_ram_bus_avalon_slave_write_pending;
  reg     [  3: 0] ext_ram_bus_byteenablen /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire    [ 31: 0] ext_ram_bus_data;
  wire    [  1: 0] ext_ram_s1_counter_load_value;
  wire             ext_ram_s1_in_a_read_cycle;
  wire             ext_ram_s1_in_a_write_cycle;
  reg     [  1: 0] ext_ram_s1_wait_counter;
  wire             ext_ram_s1_wait_counter_eq_0;
  wire             ext_ram_s1_waits_for_read;
  wire             ext_ram_s1_waits_for_write;
  wire             ext_ram_s1_with_write_latency;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 31: 0] incoming_ext_ram_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  reg              ior_n_to_the_lan91c111 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              iow_n_to_the_lan91c111 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire    [  4: 0] lan91c111_s1_counter_load_value;
  wire             lan91c111_s1_in_a_read_cycle;
  wire             lan91c111_s1_in_a_write_cycle;
  reg     [  4: 0] lan91c111_s1_wait_counter;
  wire             lan91c111_s1_wait_counter_eq_0;
  wire             lan91c111_s1_waits_for_read;
  wire             lan91c111_s1_waits_for_write;
  wire             lan91c111_s1_with_write_latency;
  reg              last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1;
  reg              last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1;
  reg              last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1;
  reg              last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1;
  reg              last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1;
  reg              last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1;
  reg              last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1;
  reg              last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1;
  wire    [ 31: 0] outgoing_ext_ram_bus_data;
  wire    [  3: 0] p1_be_n_to_the_ext_ram;
  wire    [ 19: 0] p1_ext_ram_bus_address;
  wire    [  3: 0] p1_ext_ram_bus_byteenablen;
  wire             p1_ior_n_to_the_lan91c111;
  wire             p1_iow_n_to_the_lan91c111;
  wire             p1_read_n_to_the_ext_ram;
  wire             p1_reset_to_the_lan91c111;
  wire             p1_select_n_to_the_ext_ram;
  wire    [  1: 0] p1_std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire    [  1: 0] p1_std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire             p1_write_n_to_the_ext_ram;
  reg              read_n_to_the_ext_ram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              reset_to_the_lan91c111 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              select_n_to_the_ext_ram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             std_2s60_burst_4_downstream_arbiterlock;
  wire             std_2s60_burst_4_downstream_arbiterlock2;
  wire             std_2s60_burst_4_downstream_continuerequest;
  wire             std_2s60_burst_4_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_granted_lan91c111_s1;
  wire             std_2s60_burst_4_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1;
  reg     [  1: 0] std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire             std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register_in;
  wire             std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1;
  reg     [  1: 0] std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire             std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register_in;
  wire             std_2s60_burst_4_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_4_downstream_saved_grant_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_saved_grant_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_arbiterlock;
  wire             std_2s60_burst_5_downstream_arbiterlock2;
  wire             std_2s60_burst_5_downstream_continuerequest;
  wire             std_2s60_burst_5_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_granted_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1;
  reg     [  1: 0] std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire             std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register_in;
  wire             std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1;
  reg     [  1: 0] std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire             std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register_in;
  wire             std_2s60_burst_5_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_saved_grant_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_saved_grant_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_arbiterlock;
  wire             std_2s60_burst_8_downstream_arbiterlock2;
  wire             std_2s60_burst_8_downstream_continuerequest;
  wire             std_2s60_burst_8_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_granted_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1;
  reg     [  1: 0] std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire             std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register_in;
  wire             std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1;
  reg     [  1: 0] std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire             std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register_in;
  wire             std_2s60_burst_8_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_saved_grant_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_saved_grant_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_arbiterlock;
  wire             std_2s60_burst_9_downstream_arbiterlock2;
  wire             std_2s60_burst_9_downstream_continuerequest;
  wire             std_2s60_burst_9_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_granted_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1;
  reg     [  1: 0] std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register;
  wire             std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register_in;
  wire             std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1;
  reg     [  1: 0] std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register;
  wire             std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register_in;
  wire             std_2s60_burst_9_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_saved_grant_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_saved_grant_lan91c111_s1;
  wire             time_to_write;
  wire             wait_for_ext_ram_s1_counter;
  wire             wait_for_lan91c111_s1_counter;
  reg              write_n_to_the_ext_ram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~ext_ram_bus_avalon_slave_end_xfer;
    end


  assign ext_ram_bus_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_9_downstream_qualified_request_ext_ram_s1));
  assign std_2s60_burst_4_downstream_requests_lan91c111_s1 = (0) & (std_2s60_burst_4_downstream_read | std_2s60_burst_4_downstream_write);
  //~select_n_to_the_ext_ram of type chipselect to ~p1_select_n_to_the_ext_ram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_ram <= ~0;
      else if (1)
          select_n_to_the_ext_ram <= p1_select_n_to_the_ext_ram;
    end


  assign ext_ram_bus_avalon_slave_write_pending = 0;
  //ext_ram_bus/avalon_slave read pending calc, which is an e_assign
  assign ext_ram_bus_avalon_slave_read_pending = 0;

  //ext_ram_bus_avalon_slave_arb_share_counter set values, which is an e_mux
  assign ext_ram_bus_avalon_slave_arb_share_set_values = (std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_ext_ram_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_ext_ram_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_ext_ram_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_arbitrationshare :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_arbitrationshare :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_arbitrationshare :
    (std_2s60_burst_9_downstream_granted_ext_ram_s1)? std_2s60_burst_9_downstream_arbitrationshare :
    1;

  //ext_ram_bus_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign ext_ram_bus_avalon_slave_non_bursting_master_requests = 0;

  //ext_ram_bus_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign ext_ram_bus_avalon_slave_any_bursting_master_saved_grant = std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 |
    std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 |
    std_2s60_burst_9_downstream_saved_grant_ext_ram_s1;

  //ext_ram_bus_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign ext_ram_bus_avalon_slave_arb_share_counter_next_value = ext_ram_bus_avalon_slave_firsttransfer ? (ext_ram_bus_avalon_slave_arb_share_set_values - 1) : |ext_ram_bus_avalon_slave_arb_share_counter ? (ext_ram_bus_avalon_slave_arb_share_counter - 1) : 0;

  //ext_ram_bus_avalon_slave_allgrants all slave grants, which is an e_mux
  assign ext_ram_bus_avalon_slave_allgrants = |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector |
    |ext_ram_bus_avalon_slave_grant_vector;

  //ext_ram_bus_avalon_slave_end_xfer assignment, which is an e_assign
  assign ext_ram_bus_avalon_slave_end_xfer = ~(lan91c111_s1_waits_for_read | lan91c111_s1_waits_for_write | ext_ram_s1_waits_for_read | ext_ram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave = ext_ram_bus_avalon_slave_end_xfer & (~ext_ram_bus_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ext_ram_bus_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign ext_ram_bus_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave & ext_ram_bus_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave & ~ext_ram_bus_avalon_slave_non_bursting_master_requests);

  //ext_ram_bus_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_avalon_slave_arb_share_counter <= 0;
      else if (ext_ram_bus_avalon_slave_arb_counter_enable)
          ext_ram_bus_avalon_slave_arb_share_counter <= ext_ram_bus_avalon_slave_arb_share_counter_next_value;
    end


  //ext_ram_bus_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|ext_ram_bus_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave) | (end_xfer_arb_share_counter_term_ext_ram_bus_avalon_slave & ~ext_ram_bus_avalon_slave_non_bursting_master_requests))
          ext_ram_bus_avalon_slave_slavearbiterlockenable <= |ext_ram_bus_avalon_slave_arb_share_counter_next_value;
    end


  //std_2s60_burst_4/downstream ext_ram_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_4_downstream_arbiterlock = ext_ram_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_4_downstream_continuerequest;

  //ext_ram_bus_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ext_ram_bus_avalon_slave_slavearbiterlockenable2 = |ext_ram_bus_avalon_slave_arb_share_counter_next_value;

  //std_2s60_burst_4/downstream ext_ram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_4_downstream_arbiterlock2 = ext_ram_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_4_downstream_continuerequest;

  //std_2s60_burst_5/downstream ext_ram_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_5_downstream_arbiterlock = ext_ram_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_5_downstream_continuerequest;

  //std_2s60_burst_5/downstream ext_ram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_5_downstream_arbiterlock2 = ext_ram_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_5_downstream_continuerequest;

  //std_2s60_burst_5/downstream granted lan91c111/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1 <= std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1;
    end


  //std_2s60_burst_5_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_5_downstream_continuerequest = (last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_5_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1 & 1);

  //ext_ram_bus_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ext_ram_bus_avalon_slave_any_continuerequest = std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_9_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest |
    std_2s60_burst_4_downstream_continuerequest |
    std_2s60_burst_5_downstream_continuerequest |
    std_2s60_burst_8_downstream_continuerequest;

  //std_2s60_burst_8/downstream ext_ram_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_8_downstream_arbiterlock = ext_ram_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_8_downstream_continuerequest;

  //std_2s60_burst_8/downstream ext_ram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_8_downstream_arbiterlock2 = ext_ram_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_8_downstream_continuerequest;

  //std_2s60_burst_8/downstream granted lan91c111/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1 <= std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1;
    end


  //std_2s60_burst_8_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_8_downstream_continuerequest = (last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_8_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1 & 1);

  //std_2s60_burst_9/downstream ext_ram_bus/avalon_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_9_downstream_arbiterlock = ext_ram_bus_avalon_slave_slavearbiterlockenable & std_2s60_burst_9_downstream_continuerequest;

  //std_2s60_burst_9/downstream ext_ram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_9_downstream_arbiterlock2 = ext_ram_bus_avalon_slave_slavearbiterlockenable2 & std_2s60_burst_9_downstream_continuerequest;

  //std_2s60_burst_9/downstream granted lan91c111/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1 <= std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1;
    end


  //std_2s60_burst_9_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_9_downstream_continuerequest = (last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_9_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1 & 1);

  assign std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 = std_2s60_burst_4_downstream_requests_lan91c111_s1 & ~((std_2s60_burst_4_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_4_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_4_downstream_write) | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register_in = std_2s60_burst_4_downstream_granted_lan91c111_s1 & std_2s60_burst_4_downstream_read & ~lan91c111_s1_waits_for_read;

  //shift register p1 std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register = {std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register, std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register_in};

  //std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register <= p1_std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1, which is an e_mux
  assign std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1 = std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1_shift_register[1];

  //ext_ram_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_ext_ram_bus_data <= 0;
      else if (1)
          incoming_ext_ram_bus_data <= ext_ram_bus_data;
    end


  //lan91c111_s1_with_write_latency assignment, which is an e_assign
  assign lan91c111_s1_with_write_latency = in_a_write_cycle & (std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 | std_2s60_burst_9_downstream_qualified_request_lan91c111_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (lan91c111_s1_with_write_latency)? 1 :
    (ext_ram_s1_with_write_latency)? 1 :
    (lan91c111_s1_with_write_latency)? 1 :
    (ext_ram_s1_with_write_latency)? 1 :
    (lan91c111_s1_with_write_latency)? 1 :
    (ext_ram_s1_with_write_latency)? 1 :
    (lan91c111_s1_with_write_latency)? 1 :
    (ext_ram_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_ext_ram_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_ext_ram_bus_data <= 0;
      else if (1)
          d1_outgoing_ext_ram_bus_data <= outgoing_ext_ram_bus_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else if (1)
          d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_ext_ram_bus_data tristate driver, which is an e_assign
  assign ext_ram_bus_data = (d1_in_a_write_cycle)? d1_outgoing_ext_ram_bus_data:{32{1'bz}};

  //outgoing_ext_ram_bus_data mux, which is an e_mux
  assign outgoing_ext_ram_bus_data = (std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_writedata :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_writedata :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_writedata :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_writedata :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_writedata :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_writedata :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_writedata :
    std_2s60_burst_9_downstream_writedata;

  assign std_2s60_burst_4_downstream_requests_ext_ram_s1 = (1) & (std_2s60_burst_4_downstream_read | std_2s60_burst_4_downstream_write);
  //std_2s60_burst_5/downstream granted ext_ram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1 <= std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_5_downstream_granted_slave_ext_ram_s1;
    end


  //std_2s60_burst_8/downstream granted ext_ram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1 <= std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_8_downstream_granted_slave_ext_ram_s1;
    end


  //std_2s60_burst_9/downstream granted ext_ram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1 <= std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_9_downstream_granted_slave_ext_ram_s1;
    end


  assign std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 = std_2s60_burst_4_downstream_requests_ext_ram_s1 & ~((std_2s60_burst_4_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_4_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_4_downstream_write) | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register_in = std_2s60_burst_4_downstream_granted_ext_ram_s1 & std_2s60_burst_4_downstream_read & ~ext_ram_s1_waits_for_read;

  //shift register p1 std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register = {std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register, std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register_in};

  //std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register <= p1_std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1, which is an e_mux
  assign std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1 = std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1_shift_register[1];

  //ext_ram_s1_with_write_latency assignment, which is an e_assign
  assign ext_ram_s1_with_write_latency = in_a_write_cycle & (std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 | std_2s60_burst_9_downstream_qualified_request_ext_ram_s1);

  assign std_2s60_burst_5_downstream_requests_lan91c111_s1 = (0) & (std_2s60_burst_5_downstream_read | std_2s60_burst_5_downstream_write);
  //std_2s60_burst_4/downstream granted lan91c111/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1 <= std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1;
    end


  //std_2s60_burst_4_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_4_downstream_continuerequest = (last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1 & 1) |
    (last_cycle_std_2s60_burst_4_downstream_granted_slave_lan91c111_s1 & 1) |
    (last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1 & 1);

  assign std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 = std_2s60_burst_5_downstream_requests_lan91c111_s1 & ~((std_2s60_burst_5_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_5_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_5_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register_in = std_2s60_burst_5_downstream_granted_lan91c111_s1 & std_2s60_burst_5_downstream_read & ~lan91c111_s1_waits_for_read;

  //shift register p1 std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register = {std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register, std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register_in};

  //std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register <= p1_std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1, which is an e_mux
  assign std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1 = std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1_shift_register[1];

  assign std_2s60_burst_5_downstream_requests_ext_ram_s1 = (1) & (std_2s60_burst_5_downstream_read | std_2s60_burst_5_downstream_write);
  //std_2s60_burst_4/downstream granted ext_ram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1 <= std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 ? 1 : (ext_ram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_4_downstream_granted_slave_ext_ram_s1;
    end


  assign std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 = std_2s60_burst_5_downstream_requests_ext_ram_s1 & ~((std_2s60_burst_5_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_5_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_5_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register_in = std_2s60_burst_5_downstream_granted_ext_ram_s1 & std_2s60_burst_5_downstream_read & ~ext_ram_s1_waits_for_read;

  //shift register p1 std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register = {std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register, std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register_in};

  //std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register <= p1_std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1, which is an e_mux
  assign std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1 = std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1_shift_register[1];

  assign std_2s60_burst_8_downstream_requests_lan91c111_s1 = (1) & (std_2s60_burst_8_downstream_read | std_2s60_burst_8_downstream_write);
  assign std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 = std_2s60_burst_8_downstream_requests_lan91c111_s1 & ~((std_2s60_burst_8_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_8_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_8_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register_in = std_2s60_burst_8_downstream_granted_lan91c111_s1 & std_2s60_burst_8_downstream_read & ~lan91c111_s1_waits_for_read;

  //shift register p1 std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register = {std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register, std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register_in};

  //std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register <= p1_std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1, which is an e_mux
  assign std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1 = std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1_shift_register[1];

  assign std_2s60_burst_8_downstream_requests_ext_ram_s1 = (0) & (std_2s60_burst_8_downstream_read | std_2s60_burst_8_downstream_write);
  assign std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 = std_2s60_burst_8_downstream_requests_ext_ram_s1 & ~((std_2s60_burst_8_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_8_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_8_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_9_downstream_arbiterlock);
  //std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register_in = std_2s60_burst_8_downstream_granted_ext_ram_s1 & std_2s60_burst_8_downstream_read & ~ext_ram_s1_waits_for_read;

  //shift register p1 std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register = {std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register, std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register_in};

  //std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register <= p1_std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1, which is an e_mux
  assign std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1 = std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1_shift_register[1];

  assign std_2s60_burst_9_downstream_requests_lan91c111_s1 = (1) & (std_2s60_burst_9_downstream_read | std_2s60_burst_9_downstream_write);
  assign std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 = std_2s60_burst_9_downstream_requests_lan91c111_s1 & ~((std_2s60_burst_9_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_9_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_9_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock);
  //std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register_in = std_2s60_burst_9_downstream_granted_lan91c111_s1 & std_2s60_burst_9_downstream_read & ~lan91c111_s1_waits_for_read;

  //shift register p1 std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register = {std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register, std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register_in};

  //std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register <= p1_std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1, which is an e_mux
  assign std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1 = std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1_shift_register[1];

  assign std_2s60_burst_9_downstream_requests_ext_ram_s1 = (0) & (std_2s60_burst_9_downstream_read | std_2s60_burst_9_downstream_write);
  assign std_2s60_burst_9_downstream_qualified_request_ext_ram_s1 = std_2s60_burst_9_downstream_requests_ext_ram_s1 & ~((std_2s60_burst_9_downstream_read & (ext_ram_bus_avalon_slave_write_pending | (ext_ram_bus_avalon_slave_read_pending) | (2 < std_2s60_burst_9_downstream_latency_counter))) | ((ext_ram_bus_avalon_slave_read_pending) & std_2s60_burst_9_downstream_write) | std_2s60_burst_4_downstream_arbiterlock | std_2s60_burst_5_downstream_arbiterlock | std_2s60_burst_8_downstream_arbiterlock);
  //std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register_in = std_2s60_burst_9_downstream_granted_ext_ram_s1 & std_2s60_burst_9_downstream_read & ~ext_ram_s1_waits_for_read;

  //shift register p1 std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register = {std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register, std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register_in};

  //std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register <= p1_std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1, which is an e_mux
  assign std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1 = std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1_shift_register[1];

  //allow new arb cycle for ext_ram_bus/avalon_slave, which is an e_assign
  assign ext_ram_bus_avalon_slave_allow_new_arb_cycle = ~std_2s60_burst_4_downstream_arbiterlock & ~std_2s60_burst_5_downstream_arbiterlock & ~std_2s60_burst_8_downstream_arbiterlock & ~std_2s60_burst_9_downstream_arbiterlock;

  //std_2s60_burst_9/downstream assignment into master qualified-requests vector for lan91c111/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[0] = std_2s60_burst_9_downstream_qualified_request_lan91c111_s1;

  //std_2s60_burst_9/downstream grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_9_downstream_granted_lan91c111_s1 = ext_ram_bus_avalon_slave_grant_vector[0];

  //std_2s60_burst_9/downstream saved-grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 = ext_ram_bus_avalon_slave_arb_winner[0];

  //std_2s60_burst_8/downstream assignment into master qualified-requests vector for lan91c111/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[1] = std_2s60_burst_8_downstream_qualified_request_lan91c111_s1;

  //std_2s60_burst_8/downstream grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_8_downstream_granted_lan91c111_s1 = ext_ram_bus_avalon_slave_grant_vector[1];

  //std_2s60_burst_8/downstream saved-grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 = ext_ram_bus_avalon_slave_arb_winner[1];

  //std_2s60_burst_5/downstream assignment into master qualified-requests vector for lan91c111/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[2] = std_2s60_burst_5_downstream_qualified_request_lan91c111_s1;

  //std_2s60_burst_5/downstream grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_5_downstream_granted_lan91c111_s1 = ext_ram_bus_avalon_slave_grant_vector[2];

  //std_2s60_burst_5/downstream saved-grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 = ext_ram_bus_avalon_slave_arb_winner[2];

  //std_2s60_burst_4/downstream assignment into master qualified-requests vector for lan91c111/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[3] = std_2s60_burst_4_downstream_qualified_request_lan91c111_s1;

  //std_2s60_burst_4/downstream grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_4_downstream_granted_lan91c111_s1 = ext_ram_bus_avalon_slave_grant_vector[3];

  //std_2s60_burst_4/downstream saved-grant lan91c111/s1, which is an e_assign
  assign std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 = ext_ram_bus_avalon_slave_arb_winner[3];

  //std_2s60_burst_9/downstream assignment into master qualified-requests vector for ext_ram/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[4] = std_2s60_burst_9_downstream_qualified_request_ext_ram_s1;

  //std_2s60_burst_9/downstream grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_9_downstream_granted_ext_ram_s1 = ext_ram_bus_avalon_slave_grant_vector[4];

  //std_2s60_burst_9/downstream saved-grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 = ext_ram_bus_avalon_slave_arb_winner[4];

  //std_2s60_burst_8/downstream assignment into master qualified-requests vector for ext_ram/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[5] = std_2s60_burst_8_downstream_qualified_request_ext_ram_s1;

  //std_2s60_burst_8/downstream grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_8_downstream_granted_ext_ram_s1 = ext_ram_bus_avalon_slave_grant_vector[5];

  //std_2s60_burst_8/downstream saved-grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 = ext_ram_bus_avalon_slave_arb_winner[5];

  //std_2s60_burst_5/downstream assignment into master qualified-requests vector for ext_ram/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[6] = std_2s60_burst_5_downstream_qualified_request_ext_ram_s1;

  //std_2s60_burst_5/downstream grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_5_downstream_granted_ext_ram_s1 = ext_ram_bus_avalon_slave_grant_vector[6];

  //std_2s60_burst_5/downstream saved-grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 = ext_ram_bus_avalon_slave_arb_winner[6];

  //std_2s60_burst_4/downstream assignment into master qualified-requests vector for ext_ram/s1, which is an e_assign
  assign ext_ram_bus_avalon_slave_master_qreq_vector[7] = std_2s60_burst_4_downstream_qualified_request_ext_ram_s1;

  //std_2s60_burst_4/downstream grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_4_downstream_granted_ext_ram_s1 = ext_ram_bus_avalon_slave_grant_vector[7];

  //std_2s60_burst_4/downstream saved-grant ext_ram/s1, which is an e_assign
  assign std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 = ext_ram_bus_avalon_slave_arb_winner[7];

  //ext_ram_bus/avalon_slave chosen-master double-vector, which is an e_assign
  assign ext_ram_bus_avalon_slave_chosen_master_double_vector = {ext_ram_bus_avalon_slave_master_qreq_vector, ext_ram_bus_avalon_slave_master_qreq_vector} & ({~ext_ram_bus_avalon_slave_master_qreq_vector, ~ext_ram_bus_avalon_slave_master_qreq_vector} + ext_ram_bus_avalon_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign ext_ram_bus_avalon_slave_arb_winner = (ext_ram_bus_avalon_slave_allow_new_arb_cycle & | ext_ram_bus_avalon_slave_grant_vector) ? ext_ram_bus_avalon_slave_grant_vector : ext_ram_bus_avalon_slave_saved_chosen_master_vector;

  //saved ext_ram_bus_avalon_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_avalon_slave_saved_chosen_master_vector <= 0;
      else if (ext_ram_bus_avalon_slave_allow_new_arb_cycle)
          ext_ram_bus_avalon_slave_saved_chosen_master_vector <= |ext_ram_bus_avalon_slave_grant_vector ? ext_ram_bus_avalon_slave_grant_vector : ext_ram_bus_avalon_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ext_ram_bus_avalon_slave_grant_vector = {(ext_ram_bus_avalon_slave_chosen_master_double_vector[7] | ext_ram_bus_avalon_slave_chosen_master_double_vector[15]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[6] | ext_ram_bus_avalon_slave_chosen_master_double_vector[14]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[5] | ext_ram_bus_avalon_slave_chosen_master_double_vector[13]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[4] | ext_ram_bus_avalon_slave_chosen_master_double_vector[12]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[3] | ext_ram_bus_avalon_slave_chosen_master_double_vector[11]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[2] | ext_ram_bus_avalon_slave_chosen_master_double_vector[10]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[1] | ext_ram_bus_avalon_slave_chosen_master_double_vector[9]),
    (ext_ram_bus_avalon_slave_chosen_master_double_vector[0] | ext_ram_bus_avalon_slave_chosen_master_double_vector[8])};

  //ext_ram_bus/avalon_slave chosen master rotated left, which is an e_assign
  assign ext_ram_bus_avalon_slave_chosen_master_rot_left = (ext_ram_bus_avalon_slave_arb_winner << 1) ? (ext_ram_bus_avalon_slave_arb_winner << 1) : 1;

  //ext_ram_bus/avalon_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_avalon_slave_arb_addend <= 1;
      else if (|ext_ram_bus_avalon_slave_grant_vector)
          ext_ram_bus_avalon_slave_arb_addend <= ext_ram_bus_avalon_slave_end_xfer? ext_ram_bus_avalon_slave_chosen_master_rot_left : ext_ram_bus_avalon_slave_grant_vector;
    end


  //~reset_to_the_lan91c111 of type reset_n to ~p1_reset_to_the_lan91c111, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reset_to_the_lan91c111 <= ~0;
      else if (1)
          reset_to_the_lan91c111 <= p1_reset_to_the_lan91c111;
    end


  //~p1_reset_to_the_lan91c111 assignment, which is an e_assign
  assign p1_reset_to_the_lan91c111 = ~reset_n;

  //ext_ram_bus_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign ext_ram_bus_avalon_slave_firsttransfer = ext_ram_bus_avalon_slave_begins_xfer ? ext_ram_bus_avalon_slave_unreg_firsttransfer : ext_ram_bus_avalon_slave_reg_firsttransfer;

  //ext_ram_bus_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign ext_ram_bus_avalon_slave_unreg_firsttransfer = ~(ext_ram_bus_avalon_slave_slavearbiterlockenable & ext_ram_bus_avalon_slave_any_continuerequest);

  //ext_ram_bus_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (ext_ram_bus_avalon_slave_begins_xfer)
          ext_ram_bus_avalon_slave_reg_firsttransfer <= ext_ram_bus_avalon_slave_unreg_firsttransfer;
    end


  //ext_ram_bus_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ext_ram_bus_avalon_slave_beginbursttransfer_internal = ext_ram_bus_avalon_slave_begins_xfer;

  //ext_ram_bus_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ext_ram_bus_avalon_slave_arbitration_holdoff_internal = ext_ram_bus_avalon_slave_begins_xfer & ext_ram_bus_avalon_slave_firsttransfer;

  //~ior_n_to_the_lan91c111 of type read to ~p1_ior_n_to_the_lan91c111, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ior_n_to_the_lan91c111 <= ~0;
      else if (1)
          ior_n_to_the_lan91c111 <= p1_ior_n_to_the_lan91c111;
    end


  //~p1_ior_n_to_the_lan91c111 assignment, which is an e_mux
  assign p1_ior_n_to_the_lan91c111 = ~(((std_2s60_burst_4_downstream_granted_lan91c111_s1 & std_2s60_burst_4_downstream_read) | (std_2s60_burst_5_downstream_granted_lan91c111_s1 & std_2s60_burst_5_downstream_read) | (std_2s60_burst_8_downstream_granted_lan91c111_s1 & std_2s60_burst_8_downstream_read) | (std_2s60_burst_9_downstream_granted_lan91c111_s1 & std_2s60_burst_9_downstream_read))& ~ext_ram_bus_avalon_slave_begins_xfer & (lan91c111_s1_wait_counter < 28));

  //~iow_n_to_the_lan91c111 of type write to ~p1_iow_n_to_the_lan91c111, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          iow_n_to_the_lan91c111 <= ~0;
      else if (1)
          iow_n_to_the_lan91c111 <= p1_iow_n_to_the_lan91c111;
    end


  //~ext_ram_bus_byteenablen of type byteenable to ~p1_ext_ram_bus_byteenablen, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_byteenablen <= ~0;
      else if (1)
          ext_ram_bus_byteenablen <= p1_ext_ram_bus_byteenablen;
    end


  //~p1_iow_n_to_the_lan91c111 assignment, which is an e_mux
  assign p1_iow_n_to_the_lan91c111 = ~(((std_2s60_burst_4_downstream_granted_lan91c111_s1 & std_2s60_burst_4_downstream_write) | (std_2s60_burst_5_downstream_granted_lan91c111_s1 & std_2s60_burst_5_downstream_write) | (std_2s60_burst_8_downstream_granted_lan91c111_s1 & std_2s60_burst_8_downstream_write) | (std_2s60_burst_9_downstream_granted_lan91c111_s1 & std_2s60_burst_9_downstream_write)) & ~ext_ram_bus_avalon_slave_begins_xfer & (lan91c111_s1_wait_counter >= 1) & (lan91c111_s1_wait_counter < 29));

  //ext_ram_bus_address of type address to p1_ext_ram_bus_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_bus_address <= 0;
      else if (1)
          ext_ram_bus_address <= p1_ext_ram_bus_address;
    end


  //p1_ext_ram_bus_address mux, which is an e_mux
  assign p1_ext_ram_bus_address = (std_2s60_burst_4_downstream_granted_lan91c111_s1)? {std_2s60_burst_4_downstream_nativeaddress, 2'b0} :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? {std_2s60_burst_5_downstream_nativeaddress, 2'b0} :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? {std_2s60_burst_8_downstream_nativeaddress, 2'b0} :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? {std_2s60_burst_9_downstream_nativeaddress, 2'b0} :
    (std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_address_to_slave :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_address_to_slave :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_address_to_slave :
    std_2s60_burst_9_downstream_address_to_slave;

  //d1_ext_ram_bus_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ext_ram_bus_avalon_slave_end_xfer <= 1;
      else if (1)
          d1_ext_ram_bus_avalon_slave_end_xfer <= ext_ram_bus_avalon_slave_end_xfer;
    end


  //lan91c111_s1_waits_for_read in a cycle, which is an e_mux
  assign lan91c111_s1_waits_for_read = lan91c111_s1_in_a_read_cycle & wait_for_lan91c111_s1_counter;

  //lan91c111_s1_in_a_read_cycle assignment, which is an e_assign
  assign lan91c111_s1_in_a_read_cycle = (std_2s60_burst_4_downstream_granted_lan91c111_s1 & std_2s60_burst_4_downstream_read) | (std_2s60_burst_5_downstream_granted_lan91c111_s1 & std_2s60_burst_5_downstream_read) | (std_2s60_burst_8_downstream_granted_lan91c111_s1 & std_2s60_burst_8_downstream_read) | (std_2s60_burst_9_downstream_granted_lan91c111_s1 & std_2s60_burst_9_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = lan91c111_s1_in_a_read_cycle |
    ext_ram_s1_in_a_read_cycle;

  //lan91c111_s1_waits_for_write in a cycle, which is an e_mux
  assign lan91c111_s1_waits_for_write = lan91c111_s1_in_a_write_cycle & wait_for_lan91c111_s1_counter;

  //lan91c111_s1_in_a_write_cycle assignment, which is an e_assign
  assign lan91c111_s1_in_a_write_cycle = (std_2s60_burst_4_downstream_granted_lan91c111_s1 & std_2s60_burst_4_downstream_write) | (std_2s60_burst_5_downstream_granted_lan91c111_s1 & std_2s60_burst_5_downstream_write) | (std_2s60_burst_8_downstream_granted_lan91c111_s1 & std_2s60_burst_8_downstream_write) | (std_2s60_burst_9_downstream_granted_lan91c111_s1 & std_2s60_burst_9_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = lan91c111_s1_in_a_write_cycle |
    ext_ram_s1_in_a_write_cycle;

  assign lan91c111_s1_wait_counter_eq_0 = lan91c111_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lan91c111_s1_wait_counter <= 0;
      else if (1)
          lan91c111_s1_wait_counter <= lan91c111_s1_counter_load_value;
    end


  assign lan91c111_s1_counter_load_value = ((lan91c111_s1_in_a_write_cycle & ext_ram_bus_avalon_slave_begins_xfer))? 29 :
    ((lan91c111_s1_in_a_read_cycle & ext_ram_bus_avalon_slave_begins_xfer))? 28 :
    (~lan91c111_s1_wait_counter_eq_0)? lan91c111_s1_wait_counter - 1 :
    0;

  assign wait_for_lan91c111_s1_counter = ext_ram_bus_avalon_slave_begins_xfer | ~lan91c111_s1_wait_counter_eq_0;
  //~p1_ext_ram_bus_byteenablen byte enable port mux, which is an e_mux
  assign p1_ext_ram_bus_byteenablen = ~((std_2s60_burst_4_downstream_granted_lan91c111_s1)? std_2s60_burst_4_downstream_byteenable :
    (std_2s60_burst_5_downstream_granted_lan91c111_s1)? std_2s60_burst_5_downstream_byteenable :
    (std_2s60_burst_8_downstream_granted_lan91c111_s1)? std_2s60_burst_8_downstream_byteenable :
    (std_2s60_burst_9_downstream_granted_lan91c111_s1)? std_2s60_burst_9_downstream_byteenable :
    -1);

  assign p1_select_n_to_the_ext_ram = ~(std_2s60_burst_4_downstream_granted_ext_ram_s1 | std_2s60_burst_5_downstream_granted_ext_ram_s1 | std_2s60_burst_8_downstream_granted_ext_ram_s1 | std_2s60_burst_9_downstream_granted_ext_ram_s1);
  //~read_n_to_the_ext_ram of type read to ~p1_read_n_to_the_ext_ram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_n_to_the_ext_ram <= ~0;
      else if (1)
          read_n_to_the_ext_ram <= p1_read_n_to_the_ext_ram;
    end


  //~p1_read_n_to_the_ext_ram assignment, which is an e_mux
  assign p1_read_n_to_the_ext_ram = ~(((std_2s60_burst_4_downstream_granted_ext_ram_s1 & std_2s60_burst_4_downstream_read) | (std_2s60_burst_5_downstream_granted_ext_ram_s1 & std_2s60_burst_5_downstream_read) | (std_2s60_burst_8_downstream_granted_ext_ram_s1 & std_2s60_burst_8_downstream_read) | (std_2s60_burst_9_downstream_granted_ext_ram_s1 & std_2s60_burst_9_downstream_read))& ~ext_ram_bus_avalon_slave_begins_xfer);

  //~write_n_to_the_ext_ram of type write to ~p1_write_n_to_the_ext_ram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_n_to_the_ext_ram <= ~0;
      else if (1)
          write_n_to_the_ext_ram <= p1_write_n_to_the_ext_ram;
    end


  //~be_n_to_the_ext_ram of type byteenable to ~p1_be_n_to_the_ext_ram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          be_n_to_the_ext_ram <= ~0;
      else if (1)
          be_n_to_the_ext_ram <= p1_be_n_to_the_ext_ram;
    end


  //~p1_write_n_to_the_ext_ram assignment, which is an e_mux
  assign p1_write_n_to_the_ext_ram = ~(((std_2s60_burst_4_downstream_granted_ext_ram_s1 & std_2s60_burst_4_downstream_write) | (std_2s60_burst_5_downstream_granted_ext_ram_s1 & std_2s60_burst_5_downstream_write) | (std_2s60_burst_8_downstream_granted_ext_ram_s1 & std_2s60_burst_8_downstream_write) | (std_2s60_burst_9_downstream_granted_ext_ram_s1 & std_2s60_burst_9_downstream_write)) & ~ext_ram_bus_avalon_slave_begins_xfer & (ext_ram_s1_wait_counter >= 2));

  //ext_ram_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_ram_s1_waits_for_read = ext_ram_s1_in_a_read_cycle & wait_for_ext_ram_s1_counter;

  //ext_ram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_ram_s1_in_a_read_cycle = (std_2s60_burst_4_downstream_granted_ext_ram_s1 & std_2s60_burst_4_downstream_read) | (std_2s60_burst_5_downstream_granted_ext_ram_s1 & std_2s60_burst_5_downstream_read) | (std_2s60_burst_8_downstream_granted_ext_ram_s1 & std_2s60_burst_8_downstream_read) | (std_2s60_burst_9_downstream_granted_ext_ram_s1 & std_2s60_burst_9_downstream_read);

  //ext_ram_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_ram_s1_waits_for_write = ext_ram_s1_in_a_write_cycle & wait_for_ext_ram_s1_counter;

  //ext_ram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_ram_s1_in_a_write_cycle = (std_2s60_burst_4_downstream_granted_ext_ram_s1 & std_2s60_burst_4_downstream_write) | (std_2s60_burst_5_downstream_granted_ext_ram_s1 & std_2s60_burst_5_downstream_write) | (std_2s60_burst_8_downstream_granted_ext_ram_s1 & std_2s60_burst_8_downstream_write) | (std_2s60_burst_9_downstream_granted_ext_ram_s1 & std_2s60_burst_9_downstream_write);

  assign ext_ram_s1_wait_counter_eq_0 = ext_ram_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ram_s1_wait_counter <= 0;
      else if (1)
          ext_ram_s1_wait_counter <= ext_ram_s1_counter_load_value;
    end


  assign ext_ram_s1_counter_load_value = ((ext_ram_s1_in_a_write_cycle & ext_ram_bus_avalon_slave_begins_xfer))? 3 :
    ((ext_ram_s1_in_a_read_cycle & ext_ram_bus_avalon_slave_begins_xfer))? 3 :
    (~ext_ram_s1_wait_counter_eq_0)? ext_ram_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_ram_s1_counter = ext_ram_bus_avalon_slave_begins_xfer | ~ext_ram_s1_wait_counter_eq_0;
  //~p1_be_n_to_the_ext_ram byte enable port mux, which is an e_mux
  assign p1_be_n_to_the_ext_ram = ~((std_2s60_burst_4_downstream_granted_ext_ram_s1)? std_2s60_burst_4_downstream_byteenable :
    (std_2s60_burst_5_downstream_granted_ext_ram_s1)? std_2s60_burst_5_downstream_byteenable :
    (std_2s60_burst_8_downstream_granted_ext_ram_s1)? std_2s60_burst_8_downstream_byteenable :
    (std_2s60_burst_9_downstream_granted_ext_ram_s1)? std_2s60_burst_9_downstream_byteenable :
    -1);

  //first irq irq_from_the_lan91c111 register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_irq_from_the_lan91c111 <= 0;
      else if (1)
          d1_irq_from_the_lan91c111 <= irq_from_the_lan91c111;
    end



//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lan91c111/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_4_downstream_requests_lan91c111_s1 && (std_2s60_burst_4_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_4/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_4_downstream_requests_lan91c111_s1 && (std_2s60_burst_4_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //ext_ram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_5_downstream_requests_lan91c111_s1 && (std_2s60_burst_5_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_5/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_5_downstream_requests_lan91c111_s1 && (std_2s60_burst_5_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_8/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_8_downstream_requests_lan91c111_s1 && (std_2s60_burst_8_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_8/downstream drove 0 on its 'arbitrationshare' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_8/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_8_downstream_requests_lan91c111_s1 && (std_2s60_burst_8_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_8/downstream drove 0 on its 'burstcount' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_9/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_9_downstream_requests_lan91c111_s1 && (std_2s60_burst_9_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_9/downstream drove 0 on its 'arbitrationshare' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_9/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_9_downstream_requests_lan91c111_s1 && (std_2s60_burst_9_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_9/downstream drove 0 on its 'burstcount' port while accessing slave lan91c111/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_4_downstream_granted_ext_ram_s1 + std_2s60_burst_4_downstream_granted_lan91c111_s1 + std_2s60_burst_5_downstream_granted_ext_ram_s1 + std_2s60_burst_5_downstream_granted_lan91c111_s1 + std_2s60_burst_8_downstream_granted_ext_ram_s1 + std_2s60_burst_8_downstream_granted_lan91c111_s1 + std_2s60_burst_9_downstream_granted_ext_ram_s1 + std_2s60_burst_9_downstream_granted_lan91c111_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_4_downstream_saved_grant_ext_ram_s1 + std_2s60_burst_4_downstream_saved_grant_lan91c111_s1 + std_2s60_burst_5_downstream_saved_grant_ext_ram_s1 + std_2s60_burst_5_downstream_saved_grant_lan91c111_s1 + std_2s60_burst_8_downstream_saved_grant_ext_ram_s1 + std_2s60_burst_8_downstream_saved_grant_lan91c111_s1 + std_2s60_burst_9_downstream_saved_grant_ext_ram_s1 + std_2s60_burst_9_downstream_saved_grant_lan91c111_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_bus_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module high_res_timer_s1_arbitrator (
                                      // inputs:
                                       clk,
                                       high_res_timer_s1_irq,
                                       high_res_timer_s1_readdata,
                                       reset_n,
                                       std_2s60_burst_12_downstream_address_to_slave,
                                       std_2s60_burst_12_downstream_arbitrationshare,
                                       std_2s60_burst_12_downstream_burstcount,
                                       std_2s60_burst_12_downstream_latency_counter,
                                       std_2s60_burst_12_downstream_nativeaddress,
                                       std_2s60_burst_12_downstream_read,
                                       std_2s60_burst_12_downstream_write,
                                       std_2s60_burst_12_downstream_writedata,

                                      // outputs:
                                       d1_high_res_timer_s1_end_xfer,
                                       high_res_timer_s1_address,
                                       high_res_timer_s1_chipselect,
                                       high_res_timer_s1_irq_from_sa,
                                       high_res_timer_s1_readdata_from_sa,
                                       high_res_timer_s1_reset_n,
                                       high_res_timer_s1_write_n,
                                       high_res_timer_s1_writedata,
                                       std_2s60_burst_12_downstream_granted_high_res_timer_s1,
                                       std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1,
                                       std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1,
                                       std_2s60_burst_12_downstream_requests_high_res_timer_s1
                                    )
;

  output           d1_high_res_timer_s1_end_xfer;
  output  [  2: 0] high_res_timer_s1_address;
  output           high_res_timer_s1_chipselect;
  output           high_res_timer_s1_irq_from_sa;
  output  [ 15: 0] high_res_timer_s1_readdata_from_sa;
  output           high_res_timer_s1_reset_n;
  output           high_res_timer_s1_write_n;
  output  [ 15: 0] high_res_timer_s1_writedata;
  output           std_2s60_burst_12_downstream_granted_high_res_timer_s1;
  output           std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1;
  output           std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1;
  output           std_2s60_burst_12_downstream_requests_high_res_timer_s1;
  input            clk;
  input            high_res_timer_s1_irq;
  input   [ 15: 0] high_res_timer_s1_readdata;
  input            reset_n;
  input   [  3: 0] std_2s60_burst_12_downstream_address_to_slave;
  input   [  4: 0] std_2s60_burst_12_downstream_arbitrationshare;
  input            std_2s60_burst_12_downstream_burstcount;
  input            std_2s60_burst_12_downstream_latency_counter;
  input   [  3: 0] std_2s60_burst_12_downstream_nativeaddress;
  input            std_2s60_burst_12_downstream_read;
  input            std_2s60_burst_12_downstream_write;
  input   [ 15: 0] std_2s60_burst_12_downstream_writedata;

  reg              d1_high_res_timer_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_high_res_timer_s1;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_allgrants;
  wire             high_res_timer_s1_allow_new_arb_cycle;
  wire             high_res_timer_s1_any_bursting_master_saved_grant;
  wire             high_res_timer_s1_any_continuerequest;
  wire             high_res_timer_s1_arb_counter_enable;
  reg     [  4: 0] high_res_timer_s1_arb_share_counter;
  wire    [  4: 0] high_res_timer_s1_arb_share_counter_next_value;
  wire    [  4: 0] high_res_timer_s1_arb_share_set_values;
  wire             high_res_timer_s1_beginbursttransfer_internal;
  wire             high_res_timer_s1_begins_xfer;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_end_xfer;
  wire             high_res_timer_s1_firsttransfer;
  wire             high_res_timer_s1_grant_vector;
  wire             high_res_timer_s1_in_a_read_cycle;
  wire             high_res_timer_s1_in_a_write_cycle;
  wire             high_res_timer_s1_irq_from_sa;
  wire             high_res_timer_s1_master_qreq_vector;
  wire             high_res_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  reg              high_res_timer_s1_reg_firsttransfer;
  wire             high_res_timer_s1_reset_n;
  reg              high_res_timer_s1_slavearbiterlockenable;
  wire             high_res_timer_s1_slavearbiterlockenable2;
  wire             high_res_timer_s1_unreg_firsttransfer;
  wire             high_res_timer_s1_waits_for_read;
  wire             high_res_timer_s1_waits_for_write;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             std_2s60_burst_12_downstream_arbiterlock;
  wire             std_2s60_burst_12_downstream_arbiterlock2;
  wire             std_2s60_burst_12_downstream_continuerequest;
  wire             std_2s60_burst_12_downstream_granted_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_requests_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_saved_grant_high_res_timer_s1;
  wire             wait_for_high_res_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~high_res_timer_s1_end_xfer;
    end


  assign high_res_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1));
  //assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata;

  assign std_2s60_burst_12_downstream_requests_high_res_timer_s1 = (1) & (std_2s60_burst_12_downstream_read | std_2s60_burst_12_downstream_write);
  //high_res_timer_s1_arb_share_counter set values, which is an e_mux
  assign high_res_timer_s1_arb_share_set_values = (std_2s60_burst_12_downstream_granted_high_res_timer_s1)? std_2s60_burst_12_downstream_arbitrationshare :
    1;

  //high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign high_res_timer_s1_non_bursting_master_requests = 0;

  //high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign high_res_timer_s1_any_bursting_master_saved_grant = std_2s60_burst_12_downstream_saved_grant_high_res_timer_s1;

  //high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign high_res_timer_s1_arb_share_counter_next_value = high_res_timer_s1_firsttransfer ? (high_res_timer_s1_arb_share_set_values - 1) : |high_res_timer_s1_arb_share_counter ? (high_res_timer_s1_arb_share_counter - 1) : 0;

  //high_res_timer_s1_allgrants all slave grants, which is an e_mux
  assign high_res_timer_s1_allgrants = |high_res_timer_s1_grant_vector;

  //high_res_timer_s1_end_xfer assignment, which is an e_assign
  assign high_res_timer_s1_end_xfer = ~(high_res_timer_s1_waits_for_read | high_res_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_high_res_timer_s1 = high_res_timer_s1_end_xfer & (~high_res_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign high_res_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_high_res_timer_s1 & high_res_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests);

  //high_res_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_arb_share_counter <= 0;
      else if (high_res_timer_s1_arb_counter_enable)
          high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
    end


  //high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_slavearbiterlockenable <= 0;
      else if ((|high_res_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_high_res_timer_s1) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests))
          high_res_timer_s1_slavearbiterlockenable <= |high_res_timer_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_12/downstream high_res_timer/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_12_downstream_arbiterlock = high_res_timer_s1_slavearbiterlockenable & std_2s60_burst_12_downstream_continuerequest;

  //high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign high_res_timer_s1_slavearbiterlockenable2 = |high_res_timer_s1_arb_share_counter_next_value;

  //std_2s60_burst_12/downstream high_res_timer/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_12_downstream_arbiterlock2 = high_res_timer_s1_slavearbiterlockenable2 & std_2s60_burst_12_downstream_continuerequest;

  //high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign high_res_timer_s1_any_continuerequest = 1;

  //std_2s60_burst_12_downstream_continuerequest continued request, which is an e_assign
  assign std_2s60_burst_12_downstream_continuerequest = 1;

  assign std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 = std_2s60_burst_12_downstream_requests_high_res_timer_s1 & ~((std_2s60_burst_12_downstream_read & ((std_2s60_burst_12_downstream_latency_counter != 0))));
  //local readdatavalid std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1, which is an e_mux
  assign std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1 = std_2s60_burst_12_downstream_granted_high_res_timer_s1 & std_2s60_burst_12_downstream_read & ~high_res_timer_s1_waits_for_read;

  //high_res_timer_s1_writedata mux, which is an e_mux
  assign high_res_timer_s1_writedata = std_2s60_burst_12_downstream_writedata;

  //master is always granted when requested
  assign std_2s60_burst_12_downstream_granted_high_res_timer_s1 = std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1;

  //std_2s60_burst_12/downstream saved-grant high_res_timer/s1, which is an e_assign
  assign std_2s60_burst_12_downstream_saved_grant_high_res_timer_s1 = std_2s60_burst_12_downstream_requests_high_res_timer_s1;

  //allow new arb cycle for high_res_timer/s1, which is an e_assign
  assign high_res_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign high_res_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign high_res_timer_s1_master_qreq_vector = 1;

  //high_res_timer_s1_reset_n assignment, which is an e_assign
  assign high_res_timer_s1_reset_n = reset_n;

  assign high_res_timer_s1_chipselect = std_2s60_burst_12_downstream_granted_high_res_timer_s1;
  //high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_firsttransfer = high_res_timer_s1_begins_xfer ? high_res_timer_s1_unreg_firsttransfer : high_res_timer_s1_reg_firsttransfer;

  //high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_unreg_firsttransfer = ~(high_res_timer_s1_slavearbiterlockenable & high_res_timer_s1_any_continuerequest);

  //high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_reg_firsttransfer <= 1'b1;
      else if (high_res_timer_s1_begins_xfer)
          high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
    end


  //high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign high_res_timer_s1_beginbursttransfer_internal = high_res_timer_s1_begins_xfer;

  //~high_res_timer_s1_write_n assignment, which is an e_mux
  assign high_res_timer_s1_write_n = ~(std_2s60_burst_12_downstream_granted_high_res_timer_s1 & std_2s60_burst_12_downstream_write);

  //high_res_timer_s1_address mux, which is an e_mux
  assign high_res_timer_s1_address = std_2s60_burst_12_downstream_nativeaddress;

  //d1_high_res_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_high_res_timer_s1_end_xfer <= 1;
      else if (1)
          d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end


  //high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_read = high_res_timer_s1_in_a_read_cycle & high_res_timer_s1_begins_xfer;

  //high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_read_cycle = std_2s60_burst_12_downstream_granted_high_res_timer_s1 & std_2s60_burst_12_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = high_res_timer_s1_in_a_read_cycle;

  //high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_write = high_res_timer_s1_in_a_write_cycle & 0;

  //high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_write_cycle = std_2s60_burst_12_downstream_granted_high_res_timer_s1 & std_2s60_burst_12_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = high_res_timer_s1_in_a_write_cycle;

  assign wait_for_high_res_timer_s1_counter = 0;
  //assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //high_res_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_12/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_12_downstream_requests_high_res_timer_s1 && (std_2s60_burst_12_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_12/downstream drove 0 on its 'arbitrationshare' port while accessing slave high_res_timer/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_12/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_12_downstream_requests_high_res_timer_s1 && (std_2s60_burst_12_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_12/downstream drove 0 on its 'burstcount' port while accessing slave high_res_timer/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 reset_n,
                                                 std_2s60_burst_11_downstream_address_to_slave,
                                                 std_2s60_burst_11_downstream_arbitrationshare,
                                                 std_2s60_burst_11_downstream_burstcount,
                                                 std_2s60_burst_11_downstream_latency_counter,
                                                 std_2s60_burst_11_downstream_nativeaddress,
                                                 std_2s60_burst_11_downstream_read,
                                                 std_2s60_burst_11_downstream_write,
                                                 std_2s60_burst_11_downstream_writedata,

                                                // outputs:
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata,
                                                 std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave,
                                                 std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave
                                              )
;

  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  output           std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave;
  output           std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  output           std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave;
  input            clk;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input            reset_n;
  input   [  2: 0] std_2s60_burst_11_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_11_downstream_arbitrationshare;
  input            std_2s60_burst_11_downstream_burstcount;
  input            std_2s60_burst_11_downstream_latency_counter;
  input   [  2: 0] std_2s60_burst_11_downstream_nativeaddress;
  input            std_2s60_burst_11_downstream_read;
  input            std_2s60_burst_11_downstream_write;
  input   [ 31: 0] std_2s60_burst_11_downstream_writedata;

  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg     [  3: 0] jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire    [  3: 0] jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  3: 0] jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             std_2s60_burst_11_downstream_arbiterlock;
  wire             std_2s60_burst_11_downstream_arbiterlock2;
  wire             std_2s60_burst_11_downstream_continuerequest;
  wire             std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_saved_grant_jtag_uart_avalon_jtag_slave;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave = (1) & (std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write);
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = (std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave)? std_2s60_burst_11_downstream_arbitrationshare :
    1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = 0;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = std_2s60_burst_11_downstream_saved_grant_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //std_2s60_burst_11/downstream jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_11_downstream_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & std_2s60_burst_11_downstream_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //std_2s60_burst_11/downstream jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_11_downstream_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & std_2s60_burst_11_downstream_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //std_2s60_burst_11_downstream_continuerequest continued request, which is an e_assign
  assign std_2s60_burst_11_downstream_continuerequest = 1;

  assign std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave = std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave & ~((std_2s60_burst_11_downstream_read & ((std_2s60_burst_11_downstream_latency_counter != 0))));
  //local readdatavalid std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave = std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave & std_2s60_burst_11_downstream_read & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = std_2s60_burst_11_downstream_writedata;

  //master is always granted when requested
  assign std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave = std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave;

  //std_2s60_burst_11/downstream saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign std_2s60_burst_11_downstream_saved_grant_jtag_uart_avalon_jtag_slave = std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave & std_2s60_burst_11_downstream_read);

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave & std_2s60_burst_11_downstream_write);

  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = std_2s60_burst_11_downstream_nativeaddress;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else if (1)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave & std_2s60_burst_11_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave & std_2s60_burst_11_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_11/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave && (std_2s60_burst_11_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_11/downstream drove 0 on its 'arbitrationshare' port while accessing slave jtag_uart/avalon_jtag_slave", $time);
          $stop;
        end
    end


  //std_2s60_burst_11/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave && (std_2s60_burst_11_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_11/downstream drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_ram_64_kbytes_s1_arbitrator (
                                            // inputs:
                                             clk,
                                             onchip_ram_64_kbytes_s1_readdata,
                                             reset_n,
                                             std_2s60_burst_6_downstream_address_to_slave,
                                             std_2s60_burst_6_downstream_arbitrationshare,
                                             std_2s60_burst_6_downstream_burstcount,
                                             std_2s60_burst_6_downstream_byteenable,
                                             std_2s60_burst_6_downstream_latency_counter,
                                             std_2s60_burst_6_downstream_read,
                                             std_2s60_burst_6_downstream_write,
                                             std_2s60_burst_6_downstream_writedata,
                                             std_2s60_burst_7_downstream_address_to_slave,
                                             std_2s60_burst_7_downstream_arbitrationshare,
                                             std_2s60_burst_7_downstream_burstcount,
                                             std_2s60_burst_7_downstream_byteenable,
                                             std_2s60_burst_7_downstream_latency_counter,
                                             std_2s60_burst_7_downstream_read,
                                             std_2s60_burst_7_downstream_write,
                                             std_2s60_burst_7_downstream_writedata,

                                            // outputs:
                                             d1_onchip_ram_64_kbytes_s1_end_xfer,
                                             onchip_ram_64_kbytes_s1_address,
                                             onchip_ram_64_kbytes_s1_byteenable,
                                             onchip_ram_64_kbytes_s1_chipselect,
                                             onchip_ram_64_kbytes_s1_clken,
                                             onchip_ram_64_kbytes_s1_readdata_from_sa,
                                             onchip_ram_64_kbytes_s1_write,
                                             onchip_ram_64_kbytes_s1_writedata,
                                             std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1,
                                             std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1
                                          )
;

  output           d1_onchip_ram_64_kbytes_s1_end_xfer;
  output  [ 13: 0] onchip_ram_64_kbytes_s1_address;
  output  [  3: 0] onchip_ram_64_kbytes_s1_byteenable;
  output           onchip_ram_64_kbytes_s1_chipselect;
  output           onchip_ram_64_kbytes_s1_clken;
  output  [ 31: 0] onchip_ram_64_kbytes_s1_readdata_from_sa;
  output           onchip_ram_64_kbytes_s1_write;
  output  [ 31: 0] onchip_ram_64_kbytes_s1_writedata;
  output           std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  output           std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1;
  input            clk;
  input   [ 31: 0] onchip_ram_64_kbytes_s1_readdata;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_6_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_6_downstream_arbitrationshare;
  input            std_2s60_burst_6_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_6_downstream_byteenable;
  input            std_2s60_burst_6_downstream_latency_counter;
  input            std_2s60_burst_6_downstream_read;
  input            std_2s60_burst_6_downstream_write;
  input   [ 31: 0] std_2s60_burst_6_downstream_writedata;
  input   [ 15: 0] std_2s60_burst_7_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_7_downstream_arbitrationshare;
  input            std_2s60_burst_7_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_7_downstream_byteenable;
  input            std_2s60_burst_7_downstream_latency_counter;
  input            std_2s60_burst_7_downstream_read;
  input            std_2s60_burst_7_downstream_write;
  input   [ 31: 0] std_2s60_burst_7_downstream_writedata;

  reg              d1_onchip_ram_64_kbytes_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_std_2s60_burst_6_downstream_granted_slave_onchip_ram_64_kbytes_s1;
  reg              last_cycle_std_2s60_burst_7_downstream_granted_slave_onchip_ram_64_kbytes_s1;
  wire    [ 13: 0] onchip_ram_64_kbytes_s1_address;
  wire             onchip_ram_64_kbytes_s1_allgrants;
  wire             onchip_ram_64_kbytes_s1_allow_new_arb_cycle;
  wire             onchip_ram_64_kbytes_s1_any_bursting_master_saved_grant;
  wire             onchip_ram_64_kbytes_s1_any_continuerequest;
  reg     [  1: 0] onchip_ram_64_kbytes_s1_arb_addend;
  wire             onchip_ram_64_kbytes_s1_arb_counter_enable;
  reg     [  3: 0] onchip_ram_64_kbytes_s1_arb_share_counter;
  wire    [  3: 0] onchip_ram_64_kbytes_s1_arb_share_counter_next_value;
  wire    [  3: 0] onchip_ram_64_kbytes_s1_arb_share_set_values;
  wire    [  1: 0] onchip_ram_64_kbytes_s1_arb_winner;
  wire             onchip_ram_64_kbytes_s1_arbitration_holdoff_internal;
  wire             onchip_ram_64_kbytes_s1_beginbursttransfer_internal;
  wire             onchip_ram_64_kbytes_s1_begins_xfer;
  wire    [  3: 0] onchip_ram_64_kbytes_s1_byteenable;
  wire             onchip_ram_64_kbytes_s1_chipselect;
  wire    [  3: 0] onchip_ram_64_kbytes_s1_chosen_master_double_vector;
  wire    [  1: 0] onchip_ram_64_kbytes_s1_chosen_master_rot_left;
  wire             onchip_ram_64_kbytes_s1_clken;
  wire             onchip_ram_64_kbytes_s1_end_xfer;
  wire             onchip_ram_64_kbytes_s1_firsttransfer;
  wire    [  1: 0] onchip_ram_64_kbytes_s1_grant_vector;
  wire             onchip_ram_64_kbytes_s1_in_a_read_cycle;
  wire             onchip_ram_64_kbytes_s1_in_a_write_cycle;
  wire    [  1: 0] onchip_ram_64_kbytes_s1_master_qreq_vector;
  wire             onchip_ram_64_kbytes_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_ram_64_kbytes_s1_readdata_from_sa;
  reg              onchip_ram_64_kbytes_s1_reg_firsttransfer;
  reg     [  1: 0] onchip_ram_64_kbytes_s1_saved_chosen_master_vector;
  reg              onchip_ram_64_kbytes_s1_slavearbiterlockenable;
  wire             onchip_ram_64_kbytes_s1_slavearbiterlockenable2;
  wire             onchip_ram_64_kbytes_s1_unreg_firsttransfer;
  wire             onchip_ram_64_kbytes_s1_waits_for_read;
  wire             onchip_ram_64_kbytes_s1_waits_for_write;
  wire             onchip_ram_64_kbytes_s1_write;
  wire    [ 31: 0] onchip_ram_64_kbytes_s1_writedata;
  wire             p1_std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
  wire             p1_std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
  wire    [ 15: 0] shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_6_downstream;
  wire    [ 15: 0] shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_7_downstream;
  wire             std_2s60_burst_6_downstream_arbiterlock;
  wire             std_2s60_burst_6_downstream_arbiterlock2;
  wire             std_2s60_burst_6_downstream_continuerequest;
  wire             std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  reg              std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
  wire             std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in;
  wire             std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_arbiterlock;
  wire             std_2s60_burst_7_downstream_arbiterlock2;
  wire             std_2s60_burst_7_downstream_continuerequest;
  wire             std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  reg              std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
  wire             std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in;
  wire             std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1;
  wire             wait_for_onchip_ram_64_kbytes_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~onchip_ram_64_kbytes_s1_end_xfer;
    end


  assign onchip_ram_64_kbytes_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 | std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1));
  //assign onchip_ram_64_kbytes_s1_readdata_from_sa = onchip_ram_64_kbytes_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_ram_64_kbytes_s1_readdata_from_sa = onchip_ram_64_kbytes_s1_readdata;

  assign std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1 = (1) & (std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write);
  //onchip_ram_64_kbytes_s1_arb_share_counter set values, which is an e_mux
  assign onchip_ram_64_kbytes_s1_arb_share_set_values = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_6_downstream_arbitrationshare :
    (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_7_downstream_arbitrationshare :
    (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_6_downstream_arbitrationshare :
    (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_7_downstream_arbitrationshare :
    1;

  //onchip_ram_64_kbytes_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_ram_64_kbytes_s1_non_bursting_master_requests = 0;

  //onchip_ram_64_kbytes_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_ram_64_kbytes_s1_any_bursting_master_saved_grant = std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1 |
    std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1 |
    std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1 |
    std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1;

  //onchip_ram_64_kbytes_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_ram_64_kbytes_s1_arb_share_counter_next_value = onchip_ram_64_kbytes_s1_firsttransfer ? (onchip_ram_64_kbytes_s1_arb_share_set_values - 1) : |onchip_ram_64_kbytes_s1_arb_share_counter ? (onchip_ram_64_kbytes_s1_arb_share_counter - 1) : 0;

  //onchip_ram_64_kbytes_s1_allgrants all slave grants, which is an e_mux
  assign onchip_ram_64_kbytes_s1_allgrants = |onchip_ram_64_kbytes_s1_grant_vector |
    |onchip_ram_64_kbytes_s1_grant_vector |
    |onchip_ram_64_kbytes_s1_grant_vector |
    |onchip_ram_64_kbytes_s1_grant_vector;

  //onchip_ram_64_kbytes_s1_end_xfer assignment, which is an e_assign
  assign onchip_ram_64_kbytes_s1_end_xfer = ~(onchip_ram_64_kbytes_s1_waits_for_read | onchip_ram_64_kbytes_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1 = onchip_ram_64_kbytes_s1_end_xfer & (~onchip_ram_64_kbytes_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_ram_64_kbytes_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_ram_64_kbytes_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1 & onchip_ram_64_kbytes_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1 & ~onchip_ram_64_kbytes_s1_non_bursting_master_requests);

  //onchip_ram_64_kbytes_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_ram_64_kbytes_s1_arb_share_counter <= 0;
      else if (onchip_ram_64_kbytes_s1_arb_counter_enable)
          onchip_ram_64_kbytes_s1_arb_share_counter <= onchip_ram_64_kbytes_s1_arb_share_counter_next_value;
    end


  //onchip_ram_64_kbytes_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_ram_64_kbytes_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_ram_64_kbytes_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1) | (end_xfer_arb_share_counter_term_onchip_ram_64_kbytes_s1 & ~onchip_ram_64_kbytes_s1_non_bursting_master_requests))
          onchip_ram_64_kbytes_s1_slavearbiterlockenable <= |onchip_ram_64_kbytes_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_6/downstream onchip_ram_64_kbytes/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_6_downstream_arbiterlock = onchip_ram_64_kbytes_s1_slavearbiterlockenable & std_2s60_burst_6_downstream_continuerequest;

  //onchip_ram_64_kbytes_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_ram_64_kbytes_s1_slavearbiterlockenable2 = |onchip_ram_64_kbytes_s1_arb_share_counter_next_value;

  //std_2s60_burst_6/downstream onchip_ram_64_kbytes/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_6_downstream_arbiterlock2 = onchip_ram_64_kbytes_s1_slavearbiterlockenable2 & std_2s60_burst_6_downstream_continuerequest;

  //std_2s60_burst_7/downstream onchip_ram_64_kbytes/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_7_downstream_arbiterlock = onchip_ram_64_kbytes_s1_slavearbiterlockenable & std_2s60_burst_7_downstream_continuerequest;

  //std_2s60_burst_7/downstream onchip_ram_64_kbytes/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_7_downstream_arbiterlock2 = onchip_ram_64_kbytes_s1_slavearbiterlockenable2 & std_2s60_burst_7_downstream_continuerequest;

  //std_2s60_burst_7/downstream granted onchip_ram_64_kbytes/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_7_downstream_granted_slave_onchip_ram_64_kbytes_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_7_downstream_granted_slave_onchip_ram_64_kbytes_s1 <= std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1 ? 1 : (onchip_ram_64_kbytes_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_7_downstream_granted_slave_onchip_ram_64_kbytes_s1;
    end


  //std_2s60_burst_7_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_7_downstream_continuerequest = last_cycle_std_2s60_burst_7_downstream_granted_slave_onchip_ram_64_kbytes_s1 & 1;

  //onchip_ram_64_kbytes_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_ram_64_kbytes_s1_any_continuerequest = std_2s60_burst_7_downstream_continuerequest |
    std_2s60_burst_6_downstream_continuerequest;

  assign std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 = std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1 & ~(std_2s60_burst_7_downstream_arbiterlock);
  //std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in = std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_6_downstream_read & ~onchip_ram_64_kbytes_s1_waits_for_read;

  //shift register p1 std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register = {std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register, std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in};

  //std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register <= p1_std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1, which is an e_mux
  assign std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1 = std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;

  //onchip_ram_64_kbytes_s1_writedata mux, which is an e_mux
  assign onchip_ram_64_kbytes_s1_writedata = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_6_downstream_writedata :
    std_2s60_burst_7_downstream_writedata;

  //mux onchip_ram_64_kbytes_s1_clken, which is an e_mux
  assign onchip_ram_64_kbytes_s1_clken = 1'b1;

  assign std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1 = (1) & (std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write);
  //std_2s60_burst_6/downstream granted onchip_ram_64_kbytes/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_6_downstream_granted_slave_onchip_ram_64_kbytes_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_6_downstream_granted_slave_onchip_ram_64_kbytes_s1 <= std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1 ? 1 : (onchip_ram_64_kbytes_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_6_downstream_granted_slave_onchip_ram_64_kbytes_s1;
    end


  //std_2s60_burst_6_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_6_downstream_continuerequest = last_cycle_std_2s60_burst_6_downstream_granted_slave_onchip_ram_64_kbytes_s1 & 1;

  assign std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 = std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1 & ~(std_2s60_burst_6_downstream_arbiterlock);
  //std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in = std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_7_downstream_read & ~onchip_ram_64_kbytes_s1_waits_for_read;

  //shift register p1 std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register = {std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register, std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register_in};

  //std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register <= 0;
      else if (1)
          std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register <= p1_std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;
    end


  //local readdatavalid std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1, which is an e_mux
  assign std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1 = std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1_shift_register;

  //allow new arb cycle for onchip_ram_64_kbytes/s1, which is an e_assign
  assign onchip_ram_64_kbytes_s1_allow_new_arb_cycle = ~std_2s60_burst_6_downstream_arbiterlock & ~std_2s60_burst_7_downstream_arbiterlock;

  //std_2s60_burst_7/downstream assignment into master qualified-requests vector for onchip_ram_64_kbytes/s1, which is an e_assign
  assign onchip_ram_64_kbytes_s1_master_qreq_vector[0] = std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1;

  //std_2s60_burst_7/downstream grant onchip_ram_64_kbytes/s1, which is an e_assign
  assign std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 = onchip_ram_64_kbytes_s1_grant_vector[0];

  //std_2s60_burst_7/downstream saved-grant onchip_ram_64_kbytes/s1, which is an e_assign
  assign std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1 = onchip_ram_64_kbytes_s1_arb_winner[0];

  //std_2s60_burst_6/downstream assignment into master qualified-requests vector for onchip_ram_64_kbytes/s1, which is an e_assign
  assign onchip_ram_64_kbytes_s1_master_qreq_vector[1] = std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1;

  //std_2s60_burst_6/downstream grant onchip_ram_64_kbytes/s1, which is an e_assign
  assign std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 = onchip_ram_64_kbytes_s1_grant_vector[1];

  //std_2s60_burst_6/downstream saved-grant onchip_ram_64_kbytes/s1, which is an e_assign
  assign std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1 = onchip_ram_64_kbytes_s1_arb_winner[1];

  //onchip_ram_64_kbytes/s1 chosen-master double-vector, which is an e_assign
  assign onchip_ram_64_kbytes_s1_chosen_master_double_vector = {onchip_ram_64_kbytes_s1_master_qreq_vector, onchip_ram_64_kbytes_s1_master_qreq_vector} & ({~onchip_ram_64_kbytes_s1_master_qreq_vector, ~onchip_ram_64_kbytes_s1_master_qreq_vector} + onchip_ram_64_kbytes_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_ram_64_kbytes_s1_arb_winner = (onchip_ram_64_kbytes_s1_allow_new_arb_cycle & | onchip_ram_64_kbytes_s1_grant_vector) ? onchip_ram_64_kbytes_s1_grant_vector : onchip_ram_64_kbytes_s1_saved_chosen_master_vector;

  //saved onchip_ram_64_kbytes_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_ram_64_kbytes_s1_saved_chosen_master_vector <= 0;
      else if (onchip_ram_64_kbytes_s1_allow_new_arb_cycle)
          onchip_ram_64_kbytes_s1_saved_chosen_master_vector <= |onchip_ram_64_kbytes_s1_grant_vector ? onchip_ram_64_kbytes_s1_grant_vector : onchip_ram_64_kbytes_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_ram_64_kbytes_s1_grant_vector = {(onchip_ram_64_kbytes_s1_chosen_master_double_vector[1] | onchip_ram_64_kbytes_s1_chosen_master_double_vector[3]),
    (onchip_ram_64_kbytes_s1_chosen_master_double_vector[0] | onchip_ram_64_kbytes_s1_chosen_master_double_vector[2])};

  //onchip_ram_64_kbytes/s1 chosen master rotated left, which is an e_assign
  assign onchip_ram_64_kbytes_s1_chosen_master_rot_left = (onchip_ram_64_kbytes_s1_arb_winner << 1) ? (onchip_ram_64_kbytes_s1_arb_winner << 1) : 1;

  //onchip_ram_64_kbytes/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_ram_64_kbytes_s1_arb_addend <= 1;
      else if (|onchip_ram_64_kbytes_s1_grant_vector)
          onchip_ram_64_kbytes_s1_arb_addend <= onchip_ram_64_kbytes_s1_end_xfer? onchip_ram_64_kbytes_s1_chosen_master_rot_left : onchip_ram_64_kbytes_s1_grant_vector;
    end


  assign onchip_ram_64_kbytes_s1_chipselect = std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 | std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;
  //onchip_ram_64_kbytes_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_ram_64_kbytes_s1_firsttransfer = onchip_ram_64_kbytes_s1_begins_xfer ? onchip_ram_64_kbytes_s1_unreg_firsttransfer : onchip_ram_64_kbytes_s1_reg_firsttransfer;

  //onchip_ram_64_kbytes_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_ram_64_kbytes_s1_unreg_firsttransfer = ~(onchip_ram_64_kbytes_s1_slavearbiterlockenable & onchip_ram_64_kbytes_s1_any_continuerequest);

  //onchip_ram_64_kbytes_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_ram_64_kbytes_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_ram_64_kbytes_s1_begins_xfer)
          onchip_ram_64_kbytes_s1_reg_firsttransfer <= onchip_ram_64_kbytes_s1_unreg_firsttransfer;
    end


  //onchip_ram_64_kbytes_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_ram_64_kbytes_s1_beginbursttransfer_internal = onchip_ram_64_kbytes_s1_begins_xfer;

  //onchip_ram_64_kbytes_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_ram_64_kbytes_s1_arbitration_holdoff_internal = onchip_ram_64_kbytes_s1_begins_xfer & onchip_ram_64_kbytes_s1_firsttransfer;

  //onchip_ram_64_kbytes_s1_write assignment, which is an e_mux
  assign onchip_ram_64_kbytes_s1_write = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_6_downstream_write) | (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_7_downstream_write);

  assign shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_6_downstream = std_2s60_burst_6_downstream_address_to_slave;
  //onchip_ram_64_kbytes_s1_address mux, which is an e_mux
  assign onchip_ram_64_kbytes_s1_address = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1)? (shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_6_downstream >> 2) :
    (shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_7_downstream >> 2);

  assign shifted_address_to_onchip_ram_64_kbytes_s1_from_std_2s60_burst_7_downstream = std_2s60_burst_7_downstream_address_to_slave;
  //d1_onchip_ram_64_kbytes_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_ram_64_kbytes_s1_end_xfer <= 1;
      else if (1)
          d1_onchip_ram_64_kbytes_s1_end_xfer <= onchip_ram_64_kbytes_s1_end_xfer;
    end


  //onchip_ram_64_kbytes_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_ram_64_kbytes_s1_waits_for_read = onchip_ram_64_kbytes_s1_in_a_read_cycle & 0;

  //onchip_ram_64_kbytes_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_ram_64_kbytes_s1_in_a_read_cycle = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_6_downstream_read) | (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_7_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_ram_64_kbytes_s1_in_a_read_cycle;

  //onchip_ram_64_kbytes_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_ram_64_kbytes_s1_waits_for_write = onchip_ram_64_kbytes_s1_in_a_write_cycle & 0;

  //onchip_ram_64_kbytes_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_ram_64_kbytes_s1_in_a_write_cycle = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_6_downstream_write) | (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 & std_2s60_burst_7_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_ram_64_kbytes_s1_in_a_write_cycle;

  assign wait_for_onchip_ram_64_kbytes_s1_counter = 0;
  //onchip_ram_64_kbytes_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_ram_64_kbytes_s1_byteenable = (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_6_downstream_byteenable :
    (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1)? std_2s60_burst_7_downstream_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_ram_64_kbytes/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_6/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1 && (std_2s60_burst_6_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_6/downstream drove 0 on its 'arbitrationshare' port while accessing slave onchip_ram_64_kbytes/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_6/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1 && (std_2s60_burst_6_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_6/downstream drove 0 on its 'burstcount' port while accessing slave onchip_ram_64_kbytes/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_7/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1 && (std_2s60_burst_7_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_7/downstream drove 0 on its 'arbitrationshare' port while accessing slave onchip_ram_64_kbytes/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_7/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1 && (std_2s60_burst_7_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_7/downstream drove 0 on its 'burstcount' port while accessing slave onchip_ram_64_kbytes/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 + std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_6_downstream_saved_grant_onchip_ram_64_kbytes_s1 + std_2s60_burst_7_downstream_saved_grant_onchip_ram_64_kbytes_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module reconfig_request_pio_s1_arbitrator (
                                            // inputs:
                                             clk,
                                             reconfig_request_pio_s1_readdata,
                                             reset_n,
                                             std_2s60_burst_13_downstream_address_to_slave,
                                             std_2s60_burst_13_downstream_arbitrationshare,
                                             std_2s60_burst_13_downstream_burstcount,
                                             std_2s60_burst_13_downstream_latency_counter,
                                             std_2s60_burst_13_downstream_nativeaddress,
                                             std_2s60_burst_13_downstream_read,
                                             std_2s60_burst_13_downstream_write,
                                             std_2s60_burst_13_downstream_writedata,

                                            // outputs:
                                             d1_reconfig_request_pio_s1_end_xfer,
                                             reconfig_request_pio_s1_address,
                                             reconfig_request_pio_s1_chipselect,
                                             reconfig_request_pio_s1_readdata_from_sa,
                                             reconfig_request_pio_s1_reset_n,
                                             reconfig_request_pio_s1_write_n,
                                             reconfig_request_pio_s1_writedata,
                                             std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1,
                                             std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1,
                                             std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1,
                                             std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1
                                          )
;

  output           d1_reconfig_request_pio_s1_end_xfer;
  output  [  1: 0] reconfig_request_pio_s1_address;
  output           reconfig_request_pio_s1_chipselect;
  output           reconfig_request_pio_s1_readdata_from_sa;
  output           reconfig_request_pio_s1_reset_n;
  output           reconfig_request_pio_s1_write_n;
  output           reconfig_request_pio_s1_writedata;
  output           std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1;
  output           std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1;
  output           std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1;
  output           std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1;
  input            clk;
  input            reconfig_request_pio_s1_readdata;
  input            reset_n;
  input   [  1: 0] std_2s60_burst_13_downstream_address_to_slave;
  input   [  5: 0] std_2s60_burst_13_downstream_arbitrationshare;
  input            std_2s60_burst_13_downstream_burstcount;
  input            std_2s60_burst_13_downstream_latency_counter;
  input   [  1: 0] std_2s60_burst_13_downstream_nativeaddress;
  input            std_2s60_burst_13_downstream_read;
  input            std_2s60_burst_13_downstream_write;
  input   [  7: 0] std_2s60_burst_13_downstream_writedata;

  reg              d1_reasons_to_wait;
  reg              d1_reconfig_request_pio_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_reconfig_request_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] reconfig_request_pio_s1_address;
  wire             reconfig_request_pio_s1_allgrants;
  wire             reconfig_request_pio_s1_allow_new_arb_cycle;
  wire             reconfig_request_pio_s1_any_bursting_master_saved_grant;
  wire             reconfig_request_pio_s1_any_continuerequest;
  wire             reconfig_request_pio_s1_arb_counter_enable;
  reg     [  5: 0] reconfig_request_pio_s1_arb_share_counter;
  wire    [  5: 0] reconfig_request_pio_s1_arb_share_counter_next_value;
  wire    [  5: 0] reconfig_request_pio_s1_arb_share_set_values;
  wire             reconfig_request_pio_s1_beginbursttransfer_internal;
  wire             reconfig_request_pio_s1_begins_xfer;
  wire             reconfig_request_pio_s1_chipselect;
  wire             reconfig_request_pio_s1_end_xfer;
  wire             reconfig_request_pio_s1_firsttransfer;
  wire             reconfig_request_pio_s1_grant_vector;
  wire             reconfig_request_pio_s1_in_a_read_cycle;
  wire             reconfig_request_pio_s1_in_a_write_cycle;
  wire             reconfig_request_pio_s1_master_qreq_vector;
  wire             reconfig_request_pio_s1_non_bursting_master_requests;
  wire             reconfig_request_pio_s1_readdata_from_sa;
  reg              reconfig_request_pio_s1_reg_firsttransfer;
  wire             reconfig_request_pio_s1_reset_n;
  reg              reconfig_request_pio_s1_slavearbiterlockenable;
  wire             reconfig_request_pio_s1_slavearbiterlockenable2;
  wire             reconfig_request_pio_s1_unreg_firsttransfer;
  wire             reconfig_request_pio_s1_waits_for_read;
  wire             reconfig_request_pio_s1_waits_for_write;
  wire             reconfig_request_pio_s1_write_n;
  wire             reconfig_request_pio_s1_writedata;
  wire             std_2s60_burst_13_downstream_arbiterlock;
  wire             std_2s60_burst_13_downstream_arbiterlock2;
  wire             std_2s60_burst_13_downstream_continuerequest;
  wire             std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_saved_grant_reconfig_request_pio_s1;
  wire             wait_for_reconfig_request_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~reconfig_request_pio_s1_end_xfer;
    end


  assign reconfig_request_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1));
  //assign reconfig_request_pio_s1_readdata_from_sa = reconfig_request_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign reconfig_request_pio_s1_readdata_from_sa = reconfig_request_pio_s1_readdata;

  assign std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1 = (1) & (std_2s60_burst_13_downstream_read | std_2s60_burst_13_downstream_write);
  //reconfig_request_pio_s1_arb_share_counter set values, which is an e_mux
  assign reconfig_request_pio_s1_arb_share_set_values = (std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1)? std_2s60_burst_13_downstream_arbitrationshare :
    1;

  //reconfig_request_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign reconfig_request_pio_s1_non_bursting_master_requests = 0;

  //reconfig_request_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign reconfig_request_pio_s1_any_bursting_master_saved_grant = std_2s60_burst_13_downstream_saved_grant_reconfig_request_pio_s1;

  //reconfig_request_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign reconfig_request_pio_s1_arb_share_counter_next_value = reconfig_request_pio_s1_firsttransfer ? (reconfig_request_pio_s1_arb_share_set_values - 1) : |reconfig_request_pio_s1_arb_share_counter ? (reconfig_request_pio_s1_arb_share_counter - 1) : 0;

  //reconfig_request_pio_s1_allgrants all slave grants, which is an e_mux
  assign reconfig_request_pio_s1_allgrants = |reconfig_request_pio_s1_grant_vector;

  //reconfig_request_pio_s1_end_xfer assignment, which is an e_assign
  assign reconfig_request_pio_s1_end_xfer = ~(reconfig_request_pio_s1_waits_for_read | reconfig_request_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_reconfig_request_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_reconfig_request_pio_s1 = reconfig_request_pio_s1_end_xfer & (~reconfig_request_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //reconfig_request_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign reconfig_request_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_reconfig_request_pio_s1 & reconfig_request_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_reconfig_request_pio_s1 & ~reconfig_request_pio_s1_non_bursting_master_requests);

  //reconfig_request_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reconfig_request_pio_s1_arb_share_counter <= 0;
      else if (reconfig_request_pio_s1_arb_counter_enable)
          reconfig_request_pio_s1_arb_share_counter <= reconfig_request_pio_s1_arb_share_counter_next_value;
    end


  //reconfig_request_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reconfig_request_pio_s1_slavearbiterlockenable <= 0;
      else if ((|reconfig_request_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_reconfig_request_pio_s1) | (end_xfer_arb_share_counter_term_reconfig_request_pio_s1 & ~reconfig_request_pio_s1_non_bursting_master_requests))
          reconfig_request_pio_s1_slavearbiterlockenable <= |reconfig_request_pio_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_13/downstream reconfig_request_pio/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_13_downstream_arbiterlock = reconfig_request_pio_s1_slavearbiterlockenable & std_2s60_burst_13_downstream_continuerequest;

  //reconfig_request_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign reconfig_request_pio_s1_slavearbiterlockenable2 = |reconfig_request_pio_s1_arb_share_counter_next_value;

  //std_2s60_burst_13/downstream reconfig_request_pio/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_13_downstream_arbiterlock2 = reconfig_request_pio_s1_slavearbiterlockenable2 & std_2s60_burst_13_downstream_continuerequest;

  //reconfig_request_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign reconfig_request_pio_s1_any_continuerequest = 1;

  //std_2s60_burst_13_downstream_continuerequest continued request, which is an e_assign
  assign std_2s60_burst_13_downstream_continuerequest = 1;

  assign std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 = std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1 & ~((std_2s60_burst_13_downstream_read & ((std_2s60_burst_13_downstream_latency_counter != 0))));
  //local readdatavalid std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1, which is an e_mux
  assign std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1 = std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1 & std_2s60_burst_13_downstream_read & ~reconfig_request_pio_s1_waits_for_read;

  //reconfig_request_pio_s1_writedata mux, which is an e_mux
  assign reconfig_request_pio_s1_writedata = std_2s60_burst_13_downstream_writedata;

  //master is always granted when requested
  assign std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1 = std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1;

  //std_2s60_burst_13/downstream saved-grant reconfig_request_pio/s1, which is an e_assign
  assign std_2s60_burst_13_downstream_saved_grant_reconfig_request_pio_s1 = std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1;

  //allow new arb cycle for reconfig_request_pio/s1, which is an e_assign
  assign reconfig_request_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign reconfig_request_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign reconfig_request_pio_s1_master_qreq_vector = 1;

  //reconfig_request_pio_s1_reset_n assignment, which is an e_assign
  assign reconfig_request_pio_s1_reset_n = reset_n;

  assign reconfig_request_pio_s1_chipselect = std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1;
  //reconfig_request_pio_s1_firsttransfer first transaction, which is an e_assign
  assign reconfig_request_pio_s1_firsttransfer = reconfig_request_pio_s1_begins_xfer ? reconfig_request_pio_s1_unreg_firsttransfer : reconfig_request_pio_s1_reg_firsttransfer;

  //reconfig_request_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign reconfig_request_pio_s1_unreg_firsttransfer = ~(reconfig_request_pio_s1_slavearbiterlockenable & reconfig_request_pio_s1_any_continuerequest);

  //reconfig_request_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reconfig_request_pio_s1_reg_firsttransfer <= 1'b1;
      else if (reconfig_request_pio_s1_begins_xfer)
          reconfig_request_pio_s1_reg_firsttransfer <= reconfig_request_pio_s1_unreg_firsttransfer;
    end


  //reconfig_request_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign reconfig_request_pio_s1_beginbursttransfer_internal = reconfig_request_pio_s1_begins_xfer;

  //~reconfig_request_pio_s1_write_n assignment, which is an e_mux
  assign reconfig_request_pio_s1_write_n = ~(std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1 & std_2s60_burst_13_downstream_write);

  //reconfig_request_pio_s1_address mux, which is an e_mux
  assign reconfig_request_pio_s1_address = std_2s60_burst_13_downstream_nativeaddress;

  //d1_reconfig_request_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reconfig_request_pio_s1_end_xfer <= 1;
      else if (1)
          d1_reconfig_request_pio_s1_end_xfer <= reconfig_request_pio_s1_end_xfer;
    end


  //reconfig_request_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign reconfig_request_pio_s1_waits_for_read = reconfig_request_pio_s1_in_a_read_cycle & reconfig_request_pio_s1_begins_xfer;

  //reconfig_request_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign reconfig_request_pio_s1_in_a_read_cycle = std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1 & std_2s60_burst_13_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = reconfig_request_pio_s1_in_a_read_cycle;

  //reconfig_request_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign reconfig_request_pio_s1_waits_for_write = reconfig_request_pio_s1_in_a_write_cycle & 0;

  //reconfig_request_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign reconfig_request_pio_s1_in_a_write_cycle = std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1 & std_2s60_burst_13_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = reconfig_request_pio_s1_in_a_write_cycle;

  assign wait_for_reconfig_request_pio_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //reconfig_request_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_13/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1 && (std_2s60_burst_13_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_13/downstream drove 0 on its 'arbitrationshare' port while accessing slave reconfig_request_pio/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_13/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1 && (std_2s60_burst_13_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_13/downstream drove 0 on its 'burstcount' port while accessing slave reconfig_request_pio/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_std_2s60_burst_15_downstream_to_sdram_s1_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_std_2s60_burst_16_downstream_to_sdram_s1_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sdram_s1_arbitrator (
                             // inputs:
                              clk,
                              reset_n,
                              sdram_s1_readdata,
                              sdram_s1_readdatavalid,
                              sdram_s1_waitrequest,
                              std_2s60_burst_15_downstream_address_to_slave,
                              std_2s60_burst_15_downstream_arbitrationshare,
                              std_2s60_burst_15_downstream_burstcount,
                              std_2s60_burst_15_downstream_byteenable,
                              std_2s60_burst_15_downstream_latency_counter,
                              std_2s60_burst_15_downstream_read,
                              std_2s60_burst_15_downstream_write,
                              std_2s60_burst_15_downstream_writedata,
                              std_2s60_burst_16_downstream_address_to_slave,
                              std_2s60_burst_16_downstream_arbitrationshare,
                              std_2s60_burst_16_downstream_burstcount,
                              std_2s60_burst_16_downstream_byteenable,
                              std_2s60_burst_16_downstream_latency_counter,
                              std_2s60_burst_16_downstream_read,
                              std_2s60_burst_16_downstream_write,
                              std_2s60_burst_16_downstream_writedata,

                             // outputs:
                              d1_sdram_s1_end_xfer,
                              sdram_s1_address,
                              sdram_s1_byteenable_n,
                              sdram_s1_chipselect,
                              sdram_s1_read_n,
                              sdram_s1_readdata_from_sa,
                              sdram_s1_reset_n,
                              sdram_s1_waitrequest_from_sa,
                              sdram_s1_write_n,
                              sdram_s1_writedata,
                              std_2s60_burst_15_downstream_granted_sdram_s1,
                              std_2s60_burst_15_downstream_qualified_request_sdram_s1,
                              std_2s60_burst_15_downstream_read_data_valid_sdram_s1,
                              std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register,
                              std_2s60_burst_15_downstream_requests_sdram_s1,
                              std_2s60_burst_16_downstream_granted_sdram_s1,
                              std_2s60_burst_16_downstream_qualified_request_sdram_s1,
                              std_2s60_burst_16_downstream_read_data_valid_sdram_s1,
                              std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register,
                              std_2s60_burst_16_downstream_requests_sdram_s1
                           )
;

  output           d1_sdram_s1_end_xfer;
  output  [ 21: 0] sdram_s1_address;
  output  [  3: 0] sdram_s1_byteenable_n;
  output           sdram_s1_chipselect;
  output           sdram_s1_read_n;
  output  [ 31: 0] sdram_s1_readdata_from_sa;
  output           sdram_s1_reset_n;
  output           sdram_s1_waitrequest_from_sa;
  output           sdram_s1_write_n;
  output  [ 31: 0] sdram_s1_writedata;
  output           std_2s60_burst_15_downstream_granted_sdram_s1;
  output           std_2s60_burst_15_downstream_qualified_request_sdram_s1;
  output           std_2s60_burst_15_downstream_read_data_valid_sdram_s1;
  output           std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register;
  output           std_2s60_burst_15_downstream_requests_sdram_s1;
  output           std_2s60_burst_16_downstream_granted_sdram_s1;
  output           std_2s60_burst_16_downstream_qualified_request_sdram_s1;
  output           std_2s60_burst_16_downstream_read_data_valid_sdram_s1;
  output           std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register;
  output           std_2s60_burst_16_downstream_requests_sdram_s1;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sdram_s1_readdata;
  input            sdram_s1_readdatavalid;
  input            sdram_s1_waitrequest;
  input   [ 23: 0] std_2s60_burst_15_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_15_downstream_arbitrationshare;
  input            std_2s60_burst_15_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_15_downstream_byteenable;
  input            std_2s60_burst_15_downstream_latency_counter;
  input            std_2s60_burst_15_downstream_read;
  input            std_2s60_burst_15_downstream_write;
  input   [ 31: 0] std_2s60_burst_15_downstream_writedata;
  input   [ 23: 0] std_2s60_burst_16_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_16_downstream_arbitrationshare;
  input            std_2s60_burst_16_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_16_downstream_byteenable;
  input            std_2s60_burst_16_downstream_latency_counter;
  input            std_2s60_burst_16_downstream_read;
  input            std_2s60_burst_16_downstream_write;
  input   [ 31: 0] std_2s60_burst_16_downstream_writedata;

  reg              d1_reasons_to_wait;
  reg              d1_sdram_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sdram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_std_2s60_burst_15_downstream_granted_slave_sdram_s1;
  reg              last_cycle_std_2s60_burst_16_downstream_granted_slave_sdram_s1;
  wire    [ 21: 0] sdram_s1_address;
  wire             sdram_s1_allgrants;
  wire             sdram_s1_allow_new_arb_cycle;
  wire             sdram_s1_any_bursting_master_saved_grant;
  wire             sdram_s1_any_continuerequest;
  reg     [  1: 0] sdram_s1_arb_addend;
  wire             sdram_s1_arb_counter_enable;
  reg     [  3: 0] sdram_s1_arb_share_counter;
  wire    [  3: 0] sdram_s1_arb_share_counter_next_value;
  wire    [  3: 0] sdram_s1_arb_share_set_values;
  wire    [  1: 0] sdram_s1_arb_winner;
  wire             sdram_s1_arbitration_holdoff_internal;
  wire             sdram_s1_beginbursttransfer_internal;
  wire             sdram_s1_begins_xfer;
  wire    [  3: 0] sdram_s1_byteenable_n;
  wire             sdram_s1_chipselect;
  wire    [  3: 0] sdram_s1_chosen_master_double_vector;
  wire    [  1: 0] sdram_s1_chosen_master_rot_left;
  wire             sdram_s1_end_xfer;
  wire             sdram_s1_firsttransfer;
  wire    [  1: 0] sdram_s1_grant_vector;
  wire             sdram_s1_in_a_read_cycle;
  wire             sdram_s1_in_a_write_cycle;
  wire    [  1: 0] sdram_s1_master_qreq_vector;
  wire             sdram_s1_move_on_to_next_transaction;
  wire             sdram_s1_non_bursting_master_requests;
  wire             sdram_s1_read_n;
  wire    [ 31: 0] sdram_s1_readdata_from_sa;
  wire             sdram_s1_readdatavalid_from_sa;
  reg              sdram_s1_reg_firsttransfer;
  wire             sdram_s1_reset_n;
  reg     [  1: 0] sdram_s1_saved_chosen_master_vector;
  reg              sdram_s1_slavearbiterlockenable;
  wire             sdram_s1_slavearbiterlockenable2;
  wire             sdram_s1_unreg_firsttransfer;
  wire             sdram_s1_waitrequest_from_sa;
  wire             sdram_s1_waits_for_read;
  wire             sdram_s1_waits_for_write;
  wire             sdram_s1_write_n;
  wire    [ 31: 0] sdram_s1_writedata;
  wire    [ 23: 0] shifted_address_to_sdram_s1_from_std_2s60_burst_15_downstream;
  wire    [ 23: 0] shifted_address_to_sdram_s1_from_std_2s60_burst_16_downstream;
  wire             std_2s60_burst_15_downstream_arbiterlock;
  wire             std_2s60_burst_15_downstream_arbiterlock2;
  wire             std_2s60_burst_15_downstream_continuerequest;
  wire             std_2s60_burst_15_downstream_granted_sdram_s1;
  wire             std_2s60_burst_15_downstream_qualified_request_sdram_s1;
  wire             std_2s60_burst_15_downstream_rdv_fifo_empty_sdram_s1;
  wire             std_2s60_burst_15_downstream_rdv_fifo_output_from_sdram_s1;
  wire             std_2s60_burst_15_downstream_read_data_valid_sdram_s1;
  wire             std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register;
  wire             std_2s60_burst_15_downstream_requests_sdram_s1;
  wire             std_2s60_burst_15_downstream_saved_grant_sdram_s1;
  wire             std_2s60_burst_16_downstream_arbiterlock;
  wire             std_2s60_burst_16_downstream_arbiterlock2;
  wire             std_2s60_burst_16_downstream_continuerequest;
  wire             std_2s60_burst_16_downstream_granted_sdram_s1;
  wire             std_2s60_burst_16_downstream_qualified_request_sdram_s1;
  wire             std_2s60_burst_16_downstream_rdv_fifo_empty_sdram_s1;
  wire             std_2s60_burst_16_downstream_rdv_fifo_output_from_sdram_s1;
  wire             std_2s60_burst_16_downstream_read_data_valid_sdram_s1;
  wire             std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register;
  wire             std_2s60_burst_16_downstream_requests_sdram_s1;
  wire             std_2s60_burst_16_downstream_saved_grant_sdram_s1;
  wire             wait_for_sdram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~sdram_s1_end_xfer;
    end


  assign sdram_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_15_downstream_qualified_request_sdram_s1 | std_2s60_burst_16_downstream_qualified_request_sdram_s1));
  //assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_readdata_from_sa = sdram_s1_readdata;

  assign std_2s60_burst_15_downstream_requests_sdram_s1 = (1) & (std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write);
  //assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest;

  //assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid;

  //sdram_s1_arb_share_counter set values, which is an e_mux
  assign sdram_s1_arb_share_set_values = (std_2s60_burst_15_downstream_granted_sdram_s1)? std_2s60_burst_15_downstream_arbitrationshare :
    (std_2s60_burst_16_downstream_granted_sdram_s1)? std_2s60_burst_16_downstream_arbitrationshare :
    (std_2s60_burst_15_downstream_granted_sdram_s1)? std_2s60_burst_15_downstream_arbitrationshare :
    (std_2s60_burst_16_downstream_granted_sdram_s1)? std_2s60_burst_16_downstream_arbitrationshare :
    1;

  //sdram_s1_non_bursting_master_requests mux, which is an e_mux
  assign sdram_s1_non_bursting_master_requests = 0;

  //sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sdram_s1_any_bursting_master_saved_grant = std_2s60_burst_15_downstream_saved_grant_sdram_s1 |
    std_2s60_burst_16_downstream_saved_grant_sdram_s1 |
    std_2s60_burst_15_downstream_saved_grant_sdram_s1 |
    std_2s60_burst_16_downstream_saved_grant_sdram_s1;

  //sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sdram_s1_arb_share_counter_next_value = sdram_s1_firsttransfer ? (sdram_s1_arb_share_set_values - 1) : |sdram_s1_arb_share_counter ? (sdram_s1_arb_share_counter - 1) : 0;

  //sdram_s1_allgrants all slave grants, which is an e_mux
  assign sdram_s1_allgrants = |sdram_s1_grant_vector |
    |sdram_s1_grant_vector |
    |sdram_s1_grant_vector |
    |sdram_s1_grant_vector;

  //sdram_s1_end_xfer assignment, which is an e_assign
  assign sdram_s1_end_xfer = ~(sdram_s1_waits_for_read | sdram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sdram_s1 = sdram_s1_end_xfer & (~sdram_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sdram_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sdram_s1 & sdram_s1_allgrants) | (end_xfer_arb_share_counter_term_sdram_s1 & ~sdram_s1_non_bursting_master_requests);

  //sdram_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_arb_share_counter <= 0;
      else if (sdram_s1_arb_counter_enable)
          sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
    end


  //sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_slavearbiterlockenable <= 0;
      else if ((|sdram_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sdram_s1) | (end_xfer_arb_share_counter_term_sdram_s1 & ~sdram_s1_non_bursting_master_requests))
          sdram_s1_slavearbiterlockenable <= |sdram_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_15/downstream sdram/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_15_downstream_arbiterlock = sdram_s1_slavearbiterlockenable & std_2s60_burst_15_downstream_continuerequest;

  //sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sdram_s1_slavearbiterlockenable2 = |sdram_s1_arb_share_counter_next_value;

  //std_2s60_burst_15/downstream sdram/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_15_downstream_arbiterlock2 = sdram_s1_slavearbiterlockenable2 & std_2s60_burst_15_downstream_continuerequest;

  //std_2s60_burst_16/downstream sdram/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_16_downstream_arbiterlock = sdram_s1_slavearbiterlockenable & std_2s60_burst_16_downstream_continuerequest;

  //std_2s60_burst_16/downstream sdram/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_16_downstream_arbiterlock2 = sdram_s1_slavearbiterlockenable2 & std_2s60_burst_16_downstream_continuerequest;

  //std_2s60_burst_16/downstream granted sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_16_downstream_granted_slave_sdram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_16_downstream_granted_slave_sdram_s1 <= std_2s60_burst_16_downstream_saved_grant_sdram_s1 ? 1 : (sdram_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_16_downstream_granted_slave_sdram_s1;
    end


  //std_2s60_burst_16_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_16_downstream_continuerequest = last_cycle_std_2s60_burst_16_downstream_granted_slave_sdram_s1 & 1;

  //sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sdram_s1_any_continuerequest = std_2s60_burst_16_downstream_continuerequest |
    std_2s60_burst_15_downstream_continuerequest;

  assign std_2s60_burst_15_downstream_qualified_request_sdram_s1 = std_2s60_burst_15_downstream_requests_sdram_s1 & ~((std_2s60_burst_15_downstream_read & ((std_2s60_burst_15_downstream_latency_counter != 0) | (1 < std_2s60_burst_15_downstream_latency_counter))) | std_2s60_burst_16_downstream_arbiterlock);
  //unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  assign sdram_s1_move_on_to_next_transaction = sdram_s1_readdatavalid_from_sa;

  //rdv_fifo_for_std_2s60_burst_15_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_std_2s60_burst_15_downstream_to_sdram_s1_module rdv_fifo_for_std_2s60_burst_15_downstream_to_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_15_downstream_granted_sdram_s1),
      .data_out             (std_2s60_burst_15_downstream_rdv_fifo_output_from_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (std_2s60_burst_15_downstream_rdv_fifo_empty_sdram_s1),
      .full                 (),
      .read                 (sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_s1_waits_for_read)
    );

  assign std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register = ~std_2s60_burst_15_downstream_rdv_fifo_empty_sdram_s1;
  //local readdatavalid std_2s60_burst_15_downstream_read_data_valid_sdram_s1, which is an e_mux
  assign std_2s60_burst_15_downstream_read_data_valid_sdram_s1 = (sdram_s1_readdatavalid_from_sa & std_2s60_burst_15_downstream_rdv_fifo_output_from_sdram_s1) & ~ std_2s60_burst_15_downstream_rdv_fifo_empty_sdram_s1;

  //sdram_s1_writedata mux, which is an e_mux
  assign sdram_s1_writedata = (std_2s60_burst_15_downstream_granted_sdram_s1)? std_2s60_burst_15_downstream_writedata :
    std_2s60_burst_16_downstream_writedata;

  assign std_2s60_burst_16_downstream_requests_sdram_s1 = (1) & (std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write);
  //std_2s60_burst_15/downstream granted sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_std_2s60_burst_15_downstream_granted_slave_sdram_s1 <= 0;
      else if (1)
          last_cycle_std_2s60_burst_15_downstream_granted_slave_sdram_s1 <= std_2s60_burst_15_downstream_saved_grant_sdram_s1 ? 1 : (sdram_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_std_2s60_burst_15_downstream_granted_slave_sdram_s1;
    end


  //std_2s60_burst_15_downstream_continuerequest continued request, which is an e_mux
  assign std_2s60_burst_15_downstream_continuerequest = last_cycle_std_2s60_burst_15_downstream_granted_slave_sdram_s1 & 1;

  assign std_2s60_burst_16_downstream_qualified_request_sdram_s1 = std_2s60_burst_16_downstream_requests_sdram_s1 & ~((std_2s60_burst_16_downstream_read & ((std_2s60_burst_16_downstream_latency_counter != 0) | (1 < std_2s60_burst_16_downstream_latency_counter))) | std_2s60_burst_15_downstream_arbiterlock);
  //rdv_fifo_for_std_2s60_burst_16_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_std_2s60_burst_16_downstream_to_sdram_s1_module rdv_fifo_for_std_2s60_burst_16_downstream_to_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_16_downstream_granted_sdram_s1),
      .data_out             (std_2s60_burst_16_downstream_rdv_fifo_output_from_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (std_2s60_burst_16_downstream_rdv_fifo_empty_sdram_s1),
      .full                 (),
      .read                 (sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_s1_waits_for_read)
    );

  assign std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register = ~std_2s60_burst_16_downstream_rdv_fifo_empty_sdram_s1;
  //local readdatavalid std_2s60_burst_16_downstream_read_data_valid_sdram_s1, which is an e_mux
  assign std_2s60_burst_16_downstream_read_data_valid_sdram_s1 = (sdram_s1_readdatavalid_from_sa & std_2s60_burst_16_downstream_rdv_fifo_output_from_sdram_s1) & ~ std_2s60_burst_16_downstream_rdv_fifo_empty_sdram_s1;

  //allow new arb cycle for sdram/s1, which is an e_assign
  assign sdram_s1_allow_new_arb_cycle = ~std_2s60_burst_15_downstream_arbiterlock & ~std_2s60_burst_16_downstream_arbiterlock;

  //std_2s60_burst_16/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  assign sdram_s1_master_qreq_vector[0] = std_2s60_burst_16_downstream_qualified_request_sdram_s1;

  //std_2s60_burst_16/downstream grant sdram/s1, which is an e_assign
  assign std_2s60_burst_16_downstream_granted_sdram_s1 = sdram_s1_grant_vector[0];

  //std_2s60_burst_16/downstream saved-grant sdram/s1, which is an e_assign
  assign std_2s60_burst_16_downstream_saved_grant_sdram_s1 = sdram_s1_arb_winner[0];

  //std_2s60_burst_15/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  assign sdram_s1_master_qreq_vector[1] = std_2s60_burst_15_downstream_qualified_request_sdram_s1;

  //std_2s60_burst_15/downstream grant sdram/s1, which is an e_assign
  assign std_2s60_burst_15_downstream_granted_sdram_s1 = sdram_s1_grant_vector[1];

  //std_2s60_burst_15/downstream saved-grant sdram/s1, which is an e_assign
  assign std_2s60_burst_15_downstream_saved_grant_sdram_s1 = sdram_s1_arb_winner[1];

  //sdram/s1 chosen-master double-vector, which is an e_assign
  assign sdram_s1_chosen_master_double_vector = {sdram_s1_master_qreq_vector, sdram_s1_master_qreq_vector} & ({~sdram_s1_master_qreq_vector, ~sdram_s1_master_qreq_vector} + sdram_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign sdram_s1_arb_winner = (sdram_s1_allow_new_arb_cycle & | sdram_s1_grant_vector) ? sdram_s1_grant_vector : sdram_s1_saved_chosen_master_vector;

  //saved sdram_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_saved_chosen_master_vector <= 0;
      else if (sdram_s1_allow_new_arb_cycle)
          sdram_s1_saved_chosen_master_vector <= |sdram_s1_grant_vector ? sdram_s1_grant_vector : sdram_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sdram_s1_grant_vector = {(sdram_s1_chosen_master_double_vector[1] | sdram_s1_chosen_master_double_vector[3]),
    (sdram_s1_chosen_master_double_vector[0] | sdram_s1_chosen_master_double_vector[2])};

  //sdram/s1 chosen master rotated left, which is an e_assign
  assign sdram_s1_chosen_master_rot_left = (sdram_s1_arb_winner << 1) ? (sdram_s1_arb_winner << 1) : 1;

  //sdram/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_arb_addend <= 1;
      else if (|sdram_s1_grant_vector)
          sdram_s1_arb_addend <= sdram_s1_end_xfer? sdram_s1_chosen_master_rot_left : sdram_s1_grant_vector;
    end


  //sdram_s1_reset_n assignment, which is an e_assign
  assign sdram_s1_reset_n = reset_n;

  assign sdram_s1_chipselect = std_2s60_burst_15_downstream_granted_sdram_s1 | std_2s60_burst_16_downstream_granted_sdram_s1;
  //sdram_s1_firsttransfer first transaction, which is an e_assign
  assign sdram_s1_firsttransfer = sdram_s1_begins_xfer ? sdram_s1_unreg_firsttransfer : sdram_s1_reg_firsttransfer;

  //sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sdram_s1_unreg_firsttransfer = ~(sdram_s1_slavearbiterlockenable & sdram_s1_any_continuerequest);

  //sdram_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_s1_reg_firsttransfer <= 1'b1;
      else if (sdram_s1_begins_xfer)
          sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
    end


  //sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sdram_s1_beginbursttransfer_internal = sdram_s1_begins_xfer;

  //sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sdram_s1_arbitration_holdoff_internal = sdram_s1_begins_xfer & sdram_s1_firsttransfer;

  //~sdram_s1_read_n assignment, which is an e_mux
  assign sdram_s1_read_n = ~((std_2s60_burst_15_downstream_granted_sdram_s1 & std_2s60_burst_15_downstream_read) | (std_2s60_burst_16_downstream_granted_sdram_s1 & std_2s60_burst_16_downstream_read));

  //~sdram_s1_write_n assignment, which is an e_mux
  assign sdram_s1_write_n = ~((std_2s60_burst_15_downstream_granted_sdram_s1 & std_2s60_burst_15_downstream_write) | (std_2s60_burst_16_downstream_granted_sdram_s1 & std_2s60_burst_16_downstream_write));

  assign shifted_address_to_sdram_s1_from_std_2s60_burst_15_downstream = std_2s60_burst_15_downstream_address_to_slave;
  //sdram_s1_address mux, which is an e_mux
  assign sdram_s1_address = (std_2s60_burst_15_downstream_granted_sdram_s1)? (shifted_address_to_sdram_s1_from_std_2s60_burst_15_downstream >> 2) :
    (shifted_address_to_sdram_s1_from_std_2s60_burst_16_downstream >> 2);

  assign shifted_address_to_sdram_s1_from_std_2s60_burst_16_downstream = std_2s60_burst_16_downstream_address_to_slave;
  //d1_sdram_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sdram_s1_end_xfer <= 1;
      else if (1)
          d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end


  //sdram_s1_waits_for_read in a cycle, which is an e_mux
  assign sdram_s1_waits_for_read = sdram_s1_in_a_read_cycle & sdram_s1_waitrequest_from_sa;

  //sdram_s1_in_a_read_cycle assignment, which is an e_assign
  assign sdram_s1_in_a_read_cycle = (std_2s60_burst_15_downstream_granted_sdram_s1 & std_2s60_burst_15_downstream_read) | (std_2s60_burst_16_downstream_granted_sdram_s1 & std_2s60_burst_16_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sdram_s1_in_a_read_cycle;

  //sdram_s1_waits_for_write in a cycle, which is an e_mux
  assign sdram_s1_waits_for_write = sdram_s1_in_a_write_cycle & sdram_s1_waitrequest_from_sa;

  //sdram_s1_in_a_write_cycle assignment, which is an e_assign
  assign sdram_s1_in_a_write_cycle = (std_2s60_burst_15_downstream_granted_sdram_s1 & std_2s60_burst_15_downstream_write) | (std_2s60_burst_16_downstream_granted_sdram_s1 & std_2s60_burst_16_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sdram_s1_in_a_write_cycle;

  assign wait_for_sdram_s1_counter = 0;
  //~sdram_s1_byteenable_n byte enable port mux, which is an e_mux
  assign sdram_s1_byteenable_n = ~((std_2s60_burst_15_downstream_granted_sdram_s1)? std_2s60_burst_15_downstream_byteenable :
    (std_2s60_burst_16_downstream_granted_sdram_s1)? std_2s60_burst_16_downstream_byteenable :
    -1);


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sdram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_15/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_15_downstream_requests_sdram_s1 && (std_2s60_burst_15_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_15/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_15/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_15_downstream_requests_sdram_s1 && (std_2s60_burst_15_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_15/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_16/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_16_downstream_requests_sdram_s1 && (std_2s60_burst_16_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_16/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_16/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_16_downstream_requests_sdram_s1 && (std_2s60_burst_16_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_16/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_15_downstream_granted_sdram_s1 + std_2s60_burst_16_downstream_granted_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_15_downstream_saved_grant_sdram_s1 + std_2s60_burst_16_downstream_saved_grant_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_0_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_0_upstream_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_0_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_instruction_master_address_to_slave,
                                               cpu_instruction_master_burstcount,
                                               cpu_instruction_master_latency_counter,
                                               cpu_instruction_master_read,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                               reset_n,
                                               std_2s60_burst_0_upstream_readdata,
                                               std_2s60_burst_0_upstream_readdatavalid,
                                               std_2s60_burst_0_upstream_waitrequest,

                                              // outputs:
                                               cpu_instruction_master_granted_std_2s60_burst_0_upstream,
                                               cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                               cpu_instruction_master_requests_std_2s60_burst_0_upstream,
                                               d1_std_2s60_burst_0_upstream_end_xfer,
                                               std_2s60_burst_0_upstream_address,
                                               std_2s60_burst_0_upstream_byteaddress,
                                               std_2s60_burst_0_upstream_byteenable,
                                               std_2s60_burst_0_upstream_debugaccess,
                                               std_2s60_burst_0_upstream_read,
                                               std_2s60_burst_0_upstream_readdata_from_sa,
                                               std_2s60_burst_0_upstream_waitrequest_from_sa,
                                               std_2s60_burst_0_upstream_write
                                            )
;

  output           cpu_instruction_master_granted_std_2s60_burst_0_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_0_upstream;
  output           d1_std_2s60_burst_0_upstream_end_xfer;
  output  [ 10: 0] std_2s60_burst_0_upstream_address;
  output  [ 12: 0] std_2s60_burst_0_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_0_upstream_byteenable;
  output           std_2s60_burst_0_upstream_debugaccess;
  output           std_2s60_burst_0_upstream_read;
  output  [ 31: 0] std_2s60_burst_0_upstream_readdata_from_sa;
  output           std_2s60_burst_0_upstream_waitrequest_from_sa;
  output           std_2s60_burst_0_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_0_upstream_readdata;
  input            std_2s60_burst_0_upstream_readdatavalid;
  input            std_2s60_burst_0_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_0_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_0_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_0_upstream_load_fifo;
  wire    [ 10: 0] std_2s60_burst_0_upstream_address;
  wire             std_2s60_burst_0_upstream_allgrants;
  wire             std_2s60_burst_0_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_0_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_0_upstream_any_continuerequest;
  wire             std_2s60_burst_0_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_0_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_0_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_0_upstream_arb_share_set_values;
  wire             std_2s60_burst_0_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_0_upstream_begins_xfer;
  wire             std_2s60_burst_0_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] std_2s60_burst_0_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_0_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_0_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_0_upstream_current_burst_minus_one;
  wire             std_2s60_burst_0_upstream_debugaccess;
  wire             std_2s60_burst_0_upstream_end_xfer;
  wire             std_2s60_burst_0_upstream_firsttransfer;
  wire             std_2s60_burst_0_upstream_grant_vector;
  wire             std_2s60_burst_0_upstream_in_a_read_cycle;
  wire             std_2s60_burst_0_upstream_in_a_write_cycle;
  reg              std_2s60_burst_0_upstream_load_fifo;
  wire             std_2s60_burst_0_upstream_master_qreq_vector;
  wire             std_2s60_burst_0_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_0_upstream_next_burst_count;
  wire             std_2s60_burst_0_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_0_upstream_read;
  wire    [ 31: 0] std_2s60_burst_0_upstream_readdata_from_sa;
  wire             std_2s60_burst_0_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_0_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_0_upstream_selected_burstcount;
  reg              std_2s60_burst_0_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_0_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_0_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_0_upstream_transaction_burst_count;
  wire             std_2s60_burst_0_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_0_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_0_upstream_waits_for_read;
  wire             std_2s60_burst_0_upstream_waits_for_write;
  wire             std_2s60_burst_0_upstream_write;
  wire             wait_for_std_2s60_burst_0_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_0_upstream_end_xfer;
    end


  assign std_2s60_burst_0_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream));
  //assign std_2s60_burst_0_upstream_readdata_from_sa = std_2s60_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_0_upstream_readdata_from_sa = std_2s60_burst_0_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_0_upstream = (({cpu_instruction_master_address_to_slave[25 : 11] , 11'b0} == 26'h2130800) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_0_upstream_waitrequest_from_sa = std_2s60_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_0_upstream_waitrequest_from_sa = std_2s60_burst_0_upstream_waitrequest;

  //assign std_2s60_burst_0_upstream_readdatavalid_from_sa = std_2s60_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_0_upstream_readdatavalid_from_sa = std_2s60_burst_0_upstream_readdatavalid;

  //std_2s60_burst_0_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_0_upstream_arb_share_set_values = 1;

  //std_2s60_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_0_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_0_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_0_upstream;

  //std_2s60_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_0_upstream_arb_share_counter_next_value = std_2s60_burst_0_upstream_firsttransfer ? (std_2s60_burst_0_upstream_arb_share_set_values - 1) : |std_2s60_burst_0_upstream_arb_share_counter ? (std_2s60_burst_0_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_0_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_0_upstream_allgrants = |std_2s60_burst_0_upstream_grant_vector;

  //std_2s60_burst_0_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_0_upstream_end_xfer = ~(std_2s60_burst_0_upstream_waits_for_read | std_2s60_burst_0_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream = std_2s60_burst_0_upstream_end_xfer & (~std_2s60_burst_0_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_0_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream & std_2s60_burst_0_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream & ~std_2s60_burst_0_upstream_non_bursting_master_requests);

  //std_2s60_burst_0_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_0_upstream_arb_counter_enable)
          std_2s60_burst_0_upstream_arb_share_counter <= std_2s60_burst_0_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_0_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_0_upstream & ~std_2s60_burst_0_upstream_non_bursting_master_requests))
          std_2s60_burst_0_upstream_slavearbiterlockenable <= |std_2s60_burst_0_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_0/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_0_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_0_upstream_slavearbiterlockenable2 = |std_2s60_burst_0_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_0/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_0_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_0_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream = cpu_instruction_master_requests_std_2s60_burst_0_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_0_upstream_move_on_to_next_transaction = std_2s60_burst_0_upstream_this_cycle_is_the_last_burst & std_2s60_burst_0_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_0_upstream, which is an e_mux
  assign std_2s60_burst_0_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_0_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_0_upstream_module burstcount_fifo_for_std_2s60_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_0_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_0_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_0_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_0_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read & std_2s60_burst_0_upstream_load_fifo & ~(std_2s60_burst_0_upstream_this_cycle_is_the_last_burst & std_2s60_burst_0_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_0_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_0_upstream_current_burst_minus_one = std_2s60_burst_0_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_0_upstream, which is an e_mux
  assign std_2s60_burst_0_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read) & ~std_2s60_burst_0_upstream_load_fifo))? std_2s60_burst_0_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read & std_2s60_burst_0_upstream_this_cycle_is_the_last_burst & std_2s60_burst_0_upstream_burstcount_fifo_empty))? std_2s60_burst_0_upstream_selected_burstcount :
    (std_2s60_burst_0_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_0_upstream_transaction_burst_count :
    std_2s60_burst_0_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_0_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_upstream_current_burst <= 0;
      else if (std_2s60_burst_0_upstream_readdatavalid_from_sa | (~std_2s60_burst_0_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read)))
          std_2s60_burst_0_upstream_current_burst <= std_2s60_burst_0_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_0_upstream_load_fifo = (~std_2s60_burst_0_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read) & std_2s60_burst_0_upstream_load_fifo))? 1 :
    ~std_2s60_burst_0_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read) & ~std_2s60_burst_0_upstream_load_fifo | std_2s60_burst_0_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_0_upstream_load_fifo <= p0_std_2s60_burst_0_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_0_upstream, which is an e_assign
  assign std_2s60_burst_0_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_0_upstream_current_burst_minus_one) & std_2s60_burst_0_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_0_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_0_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_0_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_0_upstream),
      .full                 (),
      .read                 (std_2s60_burst_0_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_0_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_0_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream = std_2s60_burst_0_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_0/upstream, which is an e_mux
  assign std_2s60_burst_0_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_0_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_0/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_0_upstream = cpu_instruction_master_requests_std_2s60_burst_0_upstream;

  //allow new arb cycle for std_2s60_burst_0/upstream, which is an e_assign
  assign std_2s60_burst_0_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_0_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_0_upstream_master_qreq_vector = 1;

  //std_2s60_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_0_upstream_firsttransfer = std_2s60_burst_0_upstream_begins_xfer ? std_2s60_burst_0_upstream_unreg_firsttransfer : std_2s60_burst_0_upstream_reg_firsttransfer;

  //std_2s60_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_0_upstream_unreg_firsttransfer = ~(std_2s60_burst_0_upstream_slavearbiterlockenable & std_2s60_burst_0_upstream_any_continuerequest);

  //std_2s60_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_0_upstream_begins_xfer)
          std_2s60_burst_0_upstream_reg_firsttransfer <= std_2s60_burst_0_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_0_upstream_beginbursttransfer_internal = std_2s60_burst_0_upstream_begins_xfer;

  //std_2s60_burst_0_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_0_upstream_read = cpu_instruction_master_granted_std_2s60_burst_0_upstream & cpu_instruction_master_read;

  //std_2s60_burst_0_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_0_upstream_write = 0;

  //std_2s60_burst_0_upstream_address mux, which is an e_mux
  assign std_2s60_burst_0_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_std_2s60_burst_0_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_0_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_0_upstream_end_xfer <= std_2s60_burst_0_upstream_end_xfer;
    end


  //std_2s60_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_0_upstream_waits_for_read = std_2s60_burst_0_upstream_in_a_read_cycle & std_2s60_burst_0_upstream_waitrequest_from_sa;

  //std_2s60_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_0_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_0_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_0_upstream_in_a_read_cycle;

  //std_2s60_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_0_upstream_waits_for_write = std_2s60_burst_0_upstream_in_a_write_cycle & std_2s60_burst_0_upstream_waitrequest_from_sa;

  //std_2s60_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_0_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_0_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_0_upstream_counter = 0;
  //std_2s60_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_0_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_0_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_0/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_0_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_0/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_0_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_jtag_debug_module_readdata_from_sa,
                                                 d1_cpu_jtag_debug_module_end_xfer,
                                                 reset_n,
                                                 std_2s60_burst_0_downstream_address,
                                                 std_2s60_burst_0_downstream_burstcount,
                                                 std_2s60_burst_0_downstream_byteenable,
                                                 std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module,
                                                 std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module,
                                                 std_2s60_burst_0_downstream_read,
                                                 std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module,
                                                 std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module,
                                                 std_2s60_burst_0_downstream_write,
                                                 std_2s60_burst_0_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_0_downstream_address_to_slave,
                                                 std_2s60_burst_0_downstream_latency_counter,
                                                 std_2s60_burst_0_downstream_readdata,
                                                 std_2s60_burst_0_downstream_readdatavalid,
                                                 std_2s60_burst_0_downstream_reset_n,
                                                 std_2s60_burst_0_downstream_waitrequest
                                              )
;

  output  [ 10: 0] std_2s60_burst_0_downstream_address_to_slave;
  output           std_2s60_burst_0_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_0_downstream_readdata;
  output           std_2s60_burst_0_downstream_readdatavalid;
  output           std_2s60_burst_0_downstream_reset_n;
  output           std_2s60_burst_0_downstream_waitrequest;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            reset_n;
  input   [ 10: 0] std_2s60_burst_0_downstream_address;
  input            std_2s60_burst_0_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_0_downstream_byteenable;
  input            std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module;
  input            std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  input            std_2s60_burst_0_downstream_read;
  input            std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;
  input            std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module;
  input            std_2s60_burst_0_downstream_write;
  input   [ 31: 0] std_2s60_burst_0_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_0_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_0_downstream_readdatavalid;
  wire             r_0;
  reg     [ 10: 0] std_2s60_burst_0_downstream_address_last_time;
  wire    [ 10: 0] std_2s60_burst_0_downstream_address_to_slave;
  reg              std_2s60_burst_0_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_0_downstream_byteenable_last_time;
  wire             std_2s60_burst_0_downstream_is_granted_some_slave;
  reg              std_2s60_burst_0_downstream_latency_counter;
  reg              std_2s60_burst_0_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_0_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_0_downstream_readdata;
  wire             std_2s60_burst_0_downstream_readdatavalid;
  wire             std_2s60_burst_0_downstream_reset_n;
  wire             std_2s60_burst_0_downstream_run;
  wire             std_2s60_burst_0_downstream_waitrequest;
  reg              std_2s60_burst_0_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_0_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module) & (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module | ~std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module) & ((~std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_0_downstream_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & std_2s60_burst_0_downstream_read))) & ((~std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_0_downstream_write | (1 & std_2s60_burst_0_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_0_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_0_downstream_address_to_slave = std_2s60_burst_0_downstream_address;

  //std_2s60_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_0_downstream_read_but_no_slave_selected <= std_2s60_burst_0_downstream_read & std_2s60_burst_0_downstream_run & ~std_2s60_burst_0_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_0_downstream_is_granted_some_slave = std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_0_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_0_downstream_readdatavalid = std_2s60_burst_0_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_0_downstream_readdatavalid |
    std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;

  //std_2s60_burst_0/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_0_downstream_readdata = cpu_jtag_debug_module_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_0_downstream_waitrequest = ~std_2s60_burst_0_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_0_downstream_latency_counter <= p1_std_2s60_burst_0_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_0_downstream_latency_counter = ((std_2s60_burst_0_downstream_run & std_2s60_burst_0_downstream_read))? latency_load_value :
    (std_2s60_burst_0_downstream_latency_counter)? std_2s60_burst_0_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //std_2s60_burst_0_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_0_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_0_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_address_last_time <= std_2s60_burst_0_downstream_address;
    end


  //std_2s60_burst_0/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_0_downstream_waitrequest & (std_2s60_burst_0_downstream_read | std_2s60_burst_0_downstream_write);
    end


  //std_2s60_burst_0_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_address != std_2s60_burst_0_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_0_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_burstcount_last_time <= std_2s60_burst_0_downstream_burstcount;
    end


  //std_2s60_burst_0_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_burstcount != std_2s60_burst_0_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_0_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_byteenable_last_time <= std_2s60_burst_0_downstream_byteenable;
    end


  //std_2s60_burst_0_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_byteenable != std_2s60_burst_0_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_0_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_read_last_time <= std_2s60_burst_0_downstream_read;
    end


  //std_2s60_burst_0_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_read != std_2s60_burst_0_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_0_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_write_last_time <= std_2s60_burst_0_downstream_write;
    end


  //std_2s60_burst_0_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_write != std_2s60_burst_0_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_0_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_0_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_0_downstream_writedata_last_time <= std_2s60_burst_0_downstream_writedata;
    end


  //std_2s60_burst_0_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_0_downstream_writedata != std_2s60_burst_0_downstream_writedata_last_time) & std_2s60_burst_0_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_0_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_1_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_1_upstream_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_1_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_burstcount,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_debugaccess,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                               cpu_data_master_write,
                                               cpu_data_master_writedata,
                                               reset_n,
                                               std_2s60_burst_1_upstream_readdata,
                                               std_2s60_burst_1_upstream_readdatavalid,
                                               std_2s60_burst_1_upstream_waitrequest,

                                              // outputs:
                                               cpu_data_master_granted_std_2s60_burst_1_upstream,
                                               cpu_data_master_qualified_request_std_2s60_burst_1_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                               cpu_data_master_requests_std_2s60_burst_1_upstream,
                                               d1_std_2s60_burst_1_upstream_end_xfer,
                                               std_2s60_burst_1_upstream_address,
                                               std_2s60_burst_1_upstream_burstcount,
                                               std_2s60_burst_1_upstream_byteaddress,
                                               std_2s60_burst_1_upstream_byteenable,
                                               std_2s60_burst_1_upstream_debugaccess,
                                               std_2s60_burst_1_upstream_read,
                                               std_2s60_burst_1_upstream_readdata_from_sa,
                                               std_2s60_burst_1_upstream_waitrequest_from_sa,
                                               std_2s60_burst_1_upstream_write,
                                               std_2s60_burst_1_upstream_writedata
                                            )
;

  output           cpu_data_master_granted_std_2s60_burst_1_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_1_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_1_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_1_upstream;
  output           d1_std_2s60_burst_1_upstream_end_xfer;
  output  [ 10: 0] std_2s60_burst_1_upstream_address;
  output  [  3: 0] std_2s60_burst_1_upstream_burstcount;
  output  [ 12: 0] std_2s60_burst_1_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_1_upstream_byteenable;
  output           std_2s60_burst_1_upstream_debugaccess;
  output           std_2s60_burst_1_upstream_read;
  output  [ 31: 0] std_2s60_burst_1_upstream_readdata_from_sa;
  output           std_2s60_burst_1_upstream_waitrequest_from_sa;
  output           std_2s60_burst_1_upstream_write;
  output  [ 31: 0] std_2s60_burst_1_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_1_upstream_readdata;
  input            std_2s60_burst_1_upstream_readdatavalid;
  input            std_2s60_burst_1_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_1_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_1_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_1_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_1_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_1_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_1_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_1_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_1_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_1_upstream_load_fifo;
  wire    [ 10: 0] std_2s60_burst_1_upstream_address;
  wire             std_2s60_burst_1_upstream_allgrants;
  wire             std_2s60_burst_1_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_1_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_1_upstream_any_continuerequest;
  wire             std_2s60_burst_1_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_1_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_1_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_1_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_1_upstream_bbt_burstcounter;
  wire             std_2s60_burst_1_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_1_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_1_upstream_burstcount;
  wire             std_2s60_burst_1_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] std_2s60_burst_1_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_1_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_1_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_1_upstream_current_burst_minus_one;
  wire             std_2s60_burst_1_upstream_debugaccess;
  wire             std_2s60_burst_1_upstream_end_xfer;
  wire             std_2s60_burst_1_upstream_firsttransfer;
  wire             std_2s60_burst_1_upstream_grant_vector;
  wire             std_2s60_burst_1_upstream_in_a_read_cycle;
  wire             std_2s60_burst_1_upstream_in_a_write_cycle;
  reg              std_2s60_burst_1_upstream_load_fifo;
  wire             std_2s60_burst_1_upstream_master_qreq_vector;
  wire             std_2s60_burst_1_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_1_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_1_upstream_next_burst_count;
  wire             std_2s60_burst_1_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_1_upstream_read;
  wire    [ 31: 0] std_2s60_burst_1_upstream_readdata_from_sa;
  wire             std_2s60_burst_1_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_1_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_1_upstream_selected_burstcount;
  reg              std_2s60_burst_1_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_1_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_1_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_1_upstream_transaction_burst_count;
  wire             std_2s60_burst_1_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_1_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_1_upstream_waits_for_read;
  wire             std_2s60_burst_1_upstream_waits_for_write;
  wire             std_2s60_burst_1_upstream_write;
  wire    [ 31: 0] std_2s60_burst_1_upstream_writedata;
  wire             wait_for_std_2s60_burst_1_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_1_upstream_end_xfer;
    end


  assign std_2s60_burst_1_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_1_upstream));
  //assign std_2s60_burst_1_upstream_readdata_from_sa = std_2s60_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_1_upstream_readdata_from_sa = std_2s60_burst_1_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_1_upstream = ({cpu_data_master_address_to_slave[25 : 11] , 11'b0} == 26'h2130800) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_1_upstream_waitrequest_from_sa = std_2s60_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_1_upstream_waitrequest_from_sa = std_2s60_burst_1_upstream_waitrequest;

  //assign std_2s60_burst_1_upstream_readdatavalid_from_sa = std_2s60_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_1_upstream_readdatavalid_from_sa = std_2s60_burst_1_upstream_readdatavalid;

  //std_2s60_burst_1_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_1_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_1_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_1_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_1_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_1_upstream;

  //std_2s60_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_1_upstream_arb_share_counter_next_value = std_2s60_burst_1_upstream_firsttransfer ? (std_2s60_burst_1_upstream_arb_share_set_values - 1) : |std_2s60_burst_1_upstream_arb_share_counter ? (std_2s60_burst_1_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_1_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_1_upstream_allgrants = |std_2s60_burst_1_upstream_grant_vector;

  //std_2s60_burst_1_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_1_upstream_end_xfer = ~(std_2s60_burst_1_upstream_waits_for_read | std_2s60_burst_1_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream = std_2s60_burst_1_upstream_end_xfer & (~std_2s60_burst_1_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_1_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream & std_2s60_burst_1_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream & ~std_2s60_burst_1_upstream_non_bursting_master_requests);

  //std_2s60_burst_1_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_1_upstream_arb_counter_enable)
          std_2s60_burst_1_upstream_arb_share_counter <= std_2s60_burst_1_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_1_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_1_upstream & ~std_2s60_burst_1_upstream_non_bursting_master_requests))
          std_2s60_burst_1_upstream_slavearbiterlockenable <= |std_2s60_burst_1_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_1/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_1_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_1_upstream_slavearbiterlockenable2 = |std_2s60_burst_1_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_1/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_1_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_1_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_1_upstream = cpu_data_master_requests_std_2s60_burst_1_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_1_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_1_upstream_move_on_to_next_transaction = std_2s60_burst_1_upstream_this_cycle_is_the_last_burst & std_2s60_burst_1_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_1_upstream, which is an e_mux
  assign std_2s60_burst_1_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_1_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_1_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_1_upstream_module burstcount_fifo_for_std_2s60_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_1_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_1_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_1_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_1_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read & std_2s60_burst_1_upstream_load_fifo & ~(std_2s60_burst_1_upstream_this_cycle_is_the_last_burst & std_2s60_burst_1_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_1_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_1_upstream_current_burst_minus_one = std_2s60_burst_1_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_1_upstream, which is an e_mux
  assign std_2s60_burst_1_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read) & ~std_2s60_burst_1_upstream_load_fifo))? std_2s60_burst_1_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read & std_2s60_burst_1_upstream_this_cycle_is_the_last_burst & std_2s60_burst_1_upstream_burstcount_fifo_empty))? std_2s60_burst_1_upstream_selected_burstcount :
    (std_2s60_burst_1_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_1_upstream_transaction_burst_count :
    std_2s60_burst_1_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_1_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_current_burst <= 0;
      else if (std_2s60_burst_1_upstream_readdatavalid_from_sa | (~std_2s60_burst_1_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read)))
          std_2s60_burst_1_upstream_current_burst <= std_2s60_burst_1_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_1_upstream_load_fifo = (~std_2s60_burst_1_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read) & std_2s60_burst_1_upstream_load_fifo))? 1 :
    ~std_2s60_burst_1_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read) & ~std_2s60_burst_1_upstream_load_fifo | std_2s60_burst_1_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_1_upstream_load_fifo <= p0_std_2s60_burst_1_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_1_upstream, which is an e_assign
  assign std_2s60_burst_1_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_1_upstream_current_burst_minus_one) & std_2s60_burst_1_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_1_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_1_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_1_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_1_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_1_upstream),
      .full                 (),
      .read                 (std_2s60_burst_1_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_1_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_1_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_1_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_1_upstream = std_2s60_burst_1_upstream_readdatavalid_from_sa;

  //std_2s60_burst_1_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_1_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_1/upstream, which is an e_mux
  assign std_2s60_burst_1_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_1_upstream = cpu_data_master_qualified_request_std_2s60_burst_1_upstream;

  //cpu/data_master saved-grant std_2s60_burst_1/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_1_upstream = cpu_data_master_requests_std_2s60_burst_1_upstream;

  //allow new arb cycle for std_2s60_burst_1/upstream, which is an e_assign
  assign std_2s60_burst_1_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_1_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_1_upstream_master_qreq_vector = 1;

  //std_2s60_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_1_upstream_firsttransfer = std_2s60_burst_1_upstream_begins_xfer ? std_2s60_burst_1_upstream_unreg_firsttransfer : std_2s60_burst_1_upstream_reg_firsttransfer;

  //std_2s60_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_1_upstream_unreg_firsttransfer = ~(std_2s60_burst_1_upstream_slavearbiterlockenable & std_2s60_burst_1_upstream_any_continuerequest);

  //std_2s60_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_1_upstream_begins_xfer)
          std_2s60_burst_1_upstream_reg_firsttransfer <= std_2s60_burst_1_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_1_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_1_upstream_next_bbt_burstcount = ((((std_2s60_burst_1_upstream_write) && (std_2s60_burst_1_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_1_upstream_burstcount - 1) :
    ((((std_2s60_burst_1_upstream_read) && (std_2s60_burst_1_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_1_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_1_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_1_upstream_begins_xfer)
          std_2s60_burst_1_upstream_bbt_burstcounter <= std_2s60_burst_1_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_1_upstream_beginbursttransfer_internal = std_2s60_burst_1_upstream_begins_xfer & (std_2s60_burst_1_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_1_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_1_upstream_read = cpu_data_master_granted_std_2s60_burst_1_upstream & cpu_data_master_read;

  //std_2s60_burst_1_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_1_upstream_write = cpu_data_master_granted_std_2s60_burst_1_upstream & cpu_data_master_write;

  //std_2s60_burst_1_upstream_address mux, which is an e_mux
  assign std_2s60_burst_1_upstream_address = cpu_data_master_address_to_slave;

  //d1_std_2s60_burst_1_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_1_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_1_upstream_end_xfer <= std_2s60_burst_1_upstream_end_xfer;
    end


  //std_2s60_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_1_upstream_waits_for_read = std_2s60_burst_1_upstream_in_a_read_cycle & std_2s60_burst_1_upstream_waitrequest_from_sa;

  //std_2s60_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_1_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_1_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_1_upstream_in_a_read_cycle;

  //std_2s60_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_1_upstream_waits_for_write = std_2s60_burst_1_upstream_in_a_write_cycle & std_2s60_burst_1_upstream_waitrequest_from_sa;

  //std_2s60_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_1_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_1_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_1_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_1_upstream_counter = 0;
  //std_2s60_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_1_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_1_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_1_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_1_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_1_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_1_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_1/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_1_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_1/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_1_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_jtag_debug_module_readdata_from_sa,
                                                 d1_cpu_jtag_debug_module_end_xfer,
                                                 reset_n,
                                                 std_2s60_burst_1_downstream_address,
                                                 std_2s60_burst_1_downstream_burstcount,
                                                 std_2s60_burst_1_downstream_byteenable,
                                                 std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module,
                                                 std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module,
                                                 std_2s60_burst_1_downstream_read,
                                                 std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module,
                                                 std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module,
                                                 std_2s60_burst_1_downstream_write,
                                                 std_2s60_burst_1_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_1_downstream_address_to_slave,
                                                 std_2s60_burst_1_downstream_latency_counter,
                                                 std_2s60_burst_1_downstream_readdata,
                                                 std_2s60_burst_1_downstream_readdatavalid,
                                                 std_2s60_burst_1_downstream_reset_n,
                                                 std_2s60_burst_1_downstream_waitrequest
                                              )
;

  output  [ 10: 0] std_2s60_burst_1_downstream_address_to_slave;
  output           std_2s60_burst_1_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_1_downstream_readdata;
  output           std_2s60_burst_1_downstream_readdatavalid;
  output           std_2s60_burst_1_downstream_reset_n;
  output           std_2s60_burst_1_downstream_waitrequest;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            reset_n;
  input   [ 10: 0] std_2s60_burst_1_downstream_address;
  input            std_2s60_burst_1_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_1_downstream_byteenable;
  input            std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;
  input            std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  input            std_2s60_burst_1_downstream_read;
  input            std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;
  input            std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module;
  input            std_2s60_burst_1_downstream_write;
  input   [ 31: 0] std_2s60_burst_1_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_1_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_1_downstream_readdatavalid;
  wire             r_0;
  reg     [ 10: 0] std_2s60_burst_1_downstream_address_last_time;
  wire    [ 10: 0] std_2s60_burst_1_downstream_address_to_slave;
  reg              std_2s60_burst_1_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_1_downstream_byteenable_last_time;
  wire             std_2s60_burst_1_downstream_is_granted_some_slave;
  reg              std_2s60_burst_1_downstream_latency_counter;
  reg              std_2s60_burst_1_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_1_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_1_downstream_readdata;
  wire             std_2s60_burst_1_downstream_readdatavalid;
  wire             std_2s60_burst_1_downstream_reset_n;
  wire             std_2s60_burst_1_downstream_run;
  wire             std_2s60_burst_1_downstream_waitrequest;
  reg              std_2s60_burst_1_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_1_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module) & (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module | ~std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module) & ((~std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_1_downstream_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & std_2s60_burst_1_downstream_read))) & ((~std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module | ~std_2s60_burst_1_downstream_write | (1 & std_2s60_burst_1_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_1_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_1_downstream_address_to_slave = std_2s60_burst_1_downstream_address;

  //std_2s60_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_1_downstream_read_but_no_slave_selected <= std_2s60_burst_1_downstream_read & std_2s60_burst_1_downstream_run & ~std_2s60_burst_1_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_1_downstream_is_granted_some_slave = std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_1_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_1_downstream_readdatavalid = std_2s60_burst_1_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_1_downstream_readdatavalid |
    std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;

  //std_2s60_burst_1/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_1_downstream_readdata = cpu_jtag_debug_module_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_1_downstream_waitrequest = ~std_2s60_burst_1_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_1_downstream_latency_counter <= p1_std_2s60_burst_1_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_1_downstream_latency_counter = ((std_2s60_burst_1_downstream_run & std_2s60_burst_1_downstream_read))? latency_load_value :
    (std_2s60_burst_1_downstream_latency_counter)? std_2s60_burst_1_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //std_2s60_burst_1_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_1_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_1_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_address_last_time <= std_2s60_burst_1_downstream_address;
    end


  //std_2s60_burst_1/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_1_downstream_waitrequest & (std_2s60_burst_1_downstream_read | std_2s60_burst_1_downstream_write);
    end


  //std_2s60_burst_1_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_address != std_2s60_burst_1_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_1_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_burstcount_last_time <= std_2s60_burst_1_downstream_burstcount;
    end


  //std_2s60_burst_1_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_burstcount != std_2s60_burst_1_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_1_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_byteenable_last_time <= std_2s60_burst_1_downstream_byteenable;
    end


  //std_2s60_burst_1_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_byteenable != std_2s60_burst_1_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_1_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_read_last_time <= std_2s60_burst_1_downstream_read;
    end


  //std_2s60_burst_1_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_read != std_2s60_burst_1_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_1_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_write_last_time <= std_2s60_burst_1_downstream_write;
    end


  //std_2s60_burst_1_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_write != std_2s60_burst_1_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_1_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_1_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_1_downstream_writedata_last_time <= std_2s60_burst_1_downstream_writedata;
    end


  //std_2s60_burst_1_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_1_downstream_writedata != std_2s60_burst_1_downstream_writedata_last_time) & std_2s60_burst_1_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_1_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_10_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_10_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_10_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_10_upstream_readdata,
                                                std_2s60_burst_10_upstream_readdatavalid,
                                                std_2s60_burst_10_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_10_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_10_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_10_upstream,
                                                d1_std_2s60_burst_10_upstream_end_xfer,
                                                std_2s60_burst_10_upstream_address,
                                                std_2s60_burst_10_upstream_burstcount,
                                                std_2s60_burst_10_upstream_byteaddress,
                                                std_2s60_burst_10_upstream_byteenable,
                                                std_2s60_burst_10_upstream_debugaccess,
                                                std_2s60_burst_10_upstream_read,
                                                std_2s60_burst_10_upstream_readdata_from_sa,
                                                std_2s60_burst_10_upstream_waitrequest_from_sa,
                                                std_2s60_burst_10_upstream_write,
                                                std_2s60_burst_10_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_10_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_10_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_10_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_10_upstream;
  output           d1_std_2s60_burst_10_upstream_end_xfer;
  output  [  3: 0] std_2s60_burst_10_upstream_address;
  output  [  3: 0] std_2s60_burst_10_upstream_burstcount;
  output  [  4: 0] std_2s60_burst_10_upstream_byteaddress;
  output  [  1: 0] std_2s60_burst_10_upstream_byteenable;
  output           std_2s60_burst_10_upstream_debugaccess;
  output           std_2s60_burst_10_upstream_read;
  output  [ 15: 0] std_2s60_burst_10_upstream_readdata_from_sa;
  output           std_2s60_burst_10_upstream_waitrequest_from_sa;
  output           std_2s60_burst_10_upstream_write;
  output  [ 15: 0] std_2s60_burst_10_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_10_upstream_readdata;
  input            std_2s60_burst_10_upstream_readdatavalid;
  input            std_2s60_burst_10_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_10_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_10_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_10_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_10_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_10_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_10_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_10_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_10_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_10_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_10_upstream_from_cpu_data_master;
  wire    [  3: 0] std_2s60_burst_10_upstream_address;
  wire             std_2s60_burst_10_upstream_allgrants;
  wire             std_2s60_burst_10_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_10_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_10_upstream_any_continuerequest;
  wire             std_2s60_burst_10_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_10_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_10_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_10_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_10_upstream_bbt_burstcounter;
  wire             std_2s60_burst_10_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_10_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_10_upstream_burstcount;
  wire             std_2s60_burst_10_upstream_burstcount_fifo_empty;
  wire    [  4: 0] std_2s60_burst_10_upstream_byteaddress;
  wire    [  1: 0] std_2s60_burst_10_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_10_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_10_upstream_current_burst_minus_one;
  wire             std_2s60_burst_10_upstream_debugaccess;
  wire             std_2s60_burst_10_upstream_end_xfer;
  wire             std_2s60_burst_10_upstream_firsttransfer;
  wire             std_2s60_burst_10_upstream_grant_vector;
  wire             std_2s60_burst_10_upstream_in_a_read_cycle;
  wire             std_2s60_burst_10_upstream_in_a_write_cycle;
  reg              std_2s60_burst_10_upstream_load_fifo;
  wire             std_2s60_burst_10_upstream_master_qreq_vector;
  wire             std_2s60_burst_10_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_10_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_10_upstream_next_burst_count;
  wire             std_2s60_burst_10_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_10_upstream_read;
  wire    [ 15: 0] std_2s60_burst_10_upstream_readdata_from_sa;
  wire             std_2s60_burst_10_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_10_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_10_upstream_selected_burstcount;
  reg              std_2s60_burst_10_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_10_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_10_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_10_upstream_transaction_burst_count;
  wire             std_2s60_burst_10_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_10_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_10_upstream_waits_for_read;
  wire             std_2s60_burst_10_upstream_waits_for_write;
  wire             std_2s60_burst_10_upstream_write;
  wire    [ 15: 0] std_2s60_burst_10_upstream_writedata;
  wire             wait_for_std_2s60_burst_10_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_10_upstream_end_xfer;
    end


  assign std_2s60_burst_10_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_10_upstream));
  //assign std_2s60_burst_10_upstream_readdatavalid_from_sa = std_2s60_burst_10_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_10_upstream_readdatavalid_from_sa = std_2s60_burst_10_upstream_readdatavalid;

  //assign std_2s60_burst_10_upstream_readdata_from_sa = std_2s60_burst_10_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_10_upstream_readdata_from_sa = std_2s60_burst_10_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_10_upstream = ({cpu_data_master_address_to_slave[25 : 5] , 5'b0} == 26'h2131800) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_10_upstream_waitrequest_from_sa = std_2s60_burst_10_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_10_upstream_waitrequest_from_sa = std_2s60_burst_10_upstream_waitrequest;

  //std_2s60_burst_10_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_10_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_10_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_10_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_10_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_10_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_10_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_10_upstream;

  //std_2s60_burst_10_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_10_upstream_arb_share_counter_next_value = std_2s60_burst_10_upstream_firsttransfer ? (std_2s60_burst_10_upstream_arb_share_set_values - 1) : |std_2s60_burst_10_upstream_arb_share_counter ? (std_2s60_burst_10_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_10_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_10_upstream_allgrants = |std_2s60_burst_10_upstream_grant_vector;

  //std_2s60_burst_10_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_10_upstream_end_xfer = ~(std_2s60_burst_10_upstream_waits_for_read | std_2s60_burst_10_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream = std_2s60_burst_10_upstream_end_xfer & (~std_2s60_burst_10_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_10_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_10_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream & std_2s60_burst_10_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream & ~std_2s60_burst_10_upstream_non_bursting_master_requests);

  //std_2s60_burst_10_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_10_upstream_arb_counter_enable)
          std_2s60_burst_10_upstream_arb_share_counter <= std_2s60_burst_10_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_10_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_10_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_10_upstream & ~std_2s60_burst_10_upstream_non_bursting_master_requests))
          std_2s60_burst_10_upstream_slavearbiterlockenable <= |std_2s60_burst_10_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_10/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_10_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_10_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_10_upstream_slavearbiterlockenable2 = |std_2s60_burst_10_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_10/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_10_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_10_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_10_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_10_upstream = cpu_data_master_requests_std_2s60_burst_10_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_10_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_10_upstream_move_on_to_next_transaction = std_2s60_burst_10_upstream_this_cycle_is_the_last_burst & std_2s60_burst_10_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_10_upstream, which is an e_mux
  assign std_2s60_burst_10_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_10_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_10_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_10_upstream_module burstcount_fifo_for_std_2s60_burst_10_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_10_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_10_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_10_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_10_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read & std_2s60_burst_10_upstream_load_fifo & ~(std_2s60_burst_10_upstream_this_cycle_is_the_last_burst & std_2s60_burst_10_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_10_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_10_upstream_current_burst_minus_one = std_2s60_burst_10_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_10_upstream, which is an e_mux
  assign std_2s60_burst_10_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read) & ~std_2s60_burst_10_upstream_load_fifo))? std_2s60_burst_10_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read & std_2s60_burst_10_upstream_this_cycle_is_the_last_burst & std_2s60_burst_10_upstream_burstcount_fifo_empty))? std_2s60_burst_10_upstream_selected_burstcount :
    (std_2s60_burst_10_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_10_upstream_transaction_burst_count :
    std_2s60_burst_10_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_10_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_current_burst <= 0;
      else if (std_2s60_burst_10_upstream_readdatavalid_from_sa | (~std_2s60_burst_10_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read)))
          std_2s60_burst_10_upstream_current_burst <= std_2s60_burst_10_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_10_upstream_load_fifo = (~std_2s60_burst_10_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read) & std_2s60_burst_10_upstream_load_fifo))? 1 :
    ~std_2s60_burst_10_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read) & ~std_2s60_burst_10_upstream_load_fifo | std_2s60_burst_10_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_10_upstream_load_fifo <= p0_std_2s60_burst_10_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_10_upstream, which is an e_assign
  assign std_2s60_burst_10_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_10_upstream_current_burst_minus_one) & std_2s60_burst_10_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_10_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_10_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_10_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_10_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_10_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_10_upstream),
      .full                 (),
      .read                 (std_2s60_burst_10_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_10_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_10_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_10_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_10_upstream = std_2s60_burst_10_upstream_readdatavalid_from_sa;

  //std_2s60_burst_10_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_10_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_10/upstream, which is an e_mux
  assign std_2s60_burst_10_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_10_upstream = cpu_data_master_qualified_request_std_2s60_burst_10_upstream;

  //cpu/data_master saved-grant std_2s60_burst_10/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_10_upstream = cpu_data_master_requests_std_2s60_burst_10_upstream;

  //allow new arb cycle for std_2s60_burst_10/upstream, which is an e_assign
  assign std_2s60_burst_10_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_10_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_10_upstream_master_qreq_vector = 1;

  //std_2s60_burst_10_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_10_upstream_firsttransfer = std_2s60_burst_10_upstream_begins_xfer ? std_2s60_burst_10_upstream_unreg_firsttransfer : std_2s60_burst_10_upstream_reg_firsttransfer;

  //std_2s60_burst_10_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_10_upstream_unreg_firsttransfer = ~(std_2s60_burst_10_upstream_slavearbiterlockenable & std_2s60_burst_10_upstream_any_continuerequest);

  //std_2s60_burst_10_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_10_upstream_begins_xfer)
          std_2s60_burst_10_upstream_reg_firsttransfer <= std_2s60_burst_10_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_10_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_10_upstream_next_bbt_burstcount = ((((std_2s60_burst_10_upstream_write) && (std_2s60_burst_10_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_10_upstream_burstcount - 1) :
    ((((std_2s60_burst_10_upstream_read) && (std_2s60_burst_10_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_10_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_10_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_10_upstream_begins_xfer)
          std_2s60_burst_10_upstream_bbt_burstcounter <= std_2s60_burst_10_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_10_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_10_upstream_beginbursttransfer_internal = std_2s60_burst_10_upstream_begins_xfer & (std_2s60_burst_10_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_10_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_10_upstream_read = cpu_data_master_granted_std_2s60_burst_10_upstream & cpu_data_master_read;

  //std_2s60_burst_10_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_10_upstream_write = cpu_data_master_granted_std_2s60_burst_10_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_10_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_10_upstream_address mux, which is an e_mux
  assign std_2s60_burst_10_upstream_address = shifted_address_to_std_2s60_burst_10_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_10_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_10_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_10_upstream_end_xfer <= std_2s60_burst_10_upstream_end_xfer;
    end


  //std_2s60_burst_10_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_10_upstream_waits_for_read = std_2s60_burst_10_upstream_in_a_read_cycle & std_2s60_burst_10_upstream_waitrequest_from_sa;

  //std_2s60_burst_10_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_10_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_10_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_10_upstream_in_a_read_cycle;

  //std_2s60_burst_10_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_10_upstream_waits_for_write = std_2s60_burst_10_upstream_in_a_write_cycle & std_2s60_burst_10_upstream_waitrequest_from_sa;

  //std_2s60_burst_10_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_10_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_10_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_10_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_10_upstream_counter = 0;
  //std_2s60_burst_10_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_10_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_10_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_10_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_10_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_10_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_10_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_10/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_10_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_10/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_10_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_sys_clk_timer_s1_end_xfer,
                                                  reset_n,
                                                  std_2s60_burst_10_downstream_address,
                                                  std_2s60_burst_10_downstream_burstcount,
                                                  std_2s60_burst_10_downstream_byteenable,
                                                  std_2s60_burst_10_downstream_granted_sys_clk_timer_s1,
                                                  std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1,
                                                  std_2s60_burst_10_downstream_read,
                                                  std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1,
                                                  std_2s60_burst_10_downstream_requests_sys_clk_timer_s1,
                                                  std_2s60_burst_10_downstream_write,
                                                  std_2s60_burst_10_downstream_writedata,
                                                  sys_clk_timer_s1_readdata_from_sa,

                                                 // outputs:
                                                  std_2s60_burst_10_downstream_address_to_slave,
                                                  std_2s60_burst_10_downstream_latency_counter,
                                                  std_2s60_burst_10_downstream_readdata,
                                                  std_2s60_burst_10_downstream_readdatavalid,
                                                  std_2s60_burst_10_downstream_reset_n,
                                                  std_2s60_burst_10_downstream_waitrequest
                                               )
;

  output  [  3: 0] std_2s60_burst_10_downstream_address_to_slave;
  output           std_2s60_burst_10_downstream_latency_counter;
  output  [ 15: 0] std_2s60_burst_10_downstream_readdata;
  output           std_2s60_burst_10_downstream_readdatavalid;
  output           std_2s60_burst_10_downstream_reset_n;
  output           std_2s60_burst_10_downstream_waitrequest;
  input            clk;
  input            d1_sys_clk_timer_s1_end_xfer;
  input            reset_n;
  input   [  3: 0] std_2s60_burst_10_downstream_address;
  input            std_2s60_burst_10_downstream_burstcount;
  input   [  1: 0] std_2s60_burst_10_downstream_byteenable;
  input            std_2s60_burst_10_downstream_granted_sys_clk_timer_s1;
  input            std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1;
  input            std_2s60_burst_10_downstream_read;
  input            std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1;
  input            std_2s60_burst_10_downstream_requests_sys_clk_timer_s1;
  input            std_2s60_burst_10_downstream_write;
  input   [ 15: 0] std_2s60_burst_10_downstream_writedata;
  input   [ 15: 0] sys_clk_timer_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  wire             pre_flush_std_2s60_burst_10_downstream_readdatavalid;
  wire             r_2;
  reg     [  3: 0] std_2s60_burst_10_downstream_address_last_time;
  wire    [  3: 0] std_2s60_burst_10_downstream_address_to_slave;
  reg              std_2s60_burst_10_downstream_burstcount_last_time;
  reg     [  1: 0] std_2s60_burst_10_downstream_byteenable_last_time;
  wire             std_2s60_burst_10_downstream_latency_counter;
  reg              std_2s60_burst_10_downstream_read_last_time;
  wire    [ 15: 0] std_2s60_burst_10_downstream_readdata;
  wire             std_2s60_burst_10_downstream_readdatavalid;
  wire             std_2s60_burst_10_downstream_reset_n;
  wire             std_2s60_burst_10_downstream_run;
  wire             std_2s60_burst_10_downstream_waitrequest;
  reg              std_2s60_burst_10_downstream_write_last_time;
  reg     [ 15: 0] std_2s60_burst_10_downstream_writedata_last_time;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 | ~std_2s60_burst_10_downstream_requests_sys_clk_timer_s1) & ((~std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 | ~std_2s60_burst_10_downstream_read | (1 & ~d1_sys_clk_timer_s1_end_xfer & std_2s60_burst_10_downstream_read))) & ((~std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 | ~std_2s60_burst_10_downstream_write | (1 & std_2s60_burst_10_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_10_downstream_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_10_downstream_address_to_slave = std_2s60_burst_10_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_10_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_10_downstream_readdatavalid = 0 |
    pre_flush_std_2s60_burst_10_downstream_readdatavalid |
    std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1;

  //std_2s60_burst_10/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_10_downstream_readdata = sys_clk_timer_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_10_downstream_waitrequest = ~std_2s60_burst_10_downstream_run;

  //latent max counter, which is an e_assign
  assign std_2s60_burst_10_downstream_latency_counter = 0;

  //std_2s60_burst_10_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_10_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_10_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_address_last_time <= std_2s60_burst_10_downstream_address;
    end


  //std_2s60_burst_10/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_10_downstream_waitrequest & (std_2s60_burst_10_downstream_read | std_2s60_burst_10_downstream_write);
    end


  //std_2s60_burst_10_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_address != std_2s60_burst_10_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_10_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_burstcount_last_time <= std_2s60_burst_10_downstream_burstcount;
    end


  //std_2s60_burst_10_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_burstcount != std_2s60_burst_10_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_10_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_byteenable_last_time <= std_2s60_burst_10_downstream_byteenable;
    end


  //std_2s60_burst_10_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_byteenable != std_2s60_burst_10_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_10_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_read_last_time <= std_2s60_burst_10_downstream_read;
    end


  //std_2s60_burst_10_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_read != std_2s60_burst_10_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_10_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_write_last_time <= std_2s60_burst_10_downstream_write;
    end


  //std_2s60_burst_10_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_write != std_2s60_burst_10_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_10_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_10_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_10_downstream_writedata_last_time <= std_2s60_burst_10_downstream_writedata;
    end


  //std_2s60_burst_10_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_10_downstream_writedata != std_2s60_burst_10_downstream_writedata_last_time) & std_2s60_burst_10_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_10_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_11_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_11_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_11_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_11_upstream_readdata,
                                                std_2s60_burst_11_upstream_readdatavalid,
                                                std_2s60_burst_11_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_11_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_11_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_11_upstream,
                                                d1_std_2s60_burst_11_upstream_end_xfer,
                                                std_2s60_burst_11_upstream_address,
                                                std_2s60_burst_11_upstream_burstcount,
                                                std_2s60_burst_11_upstream_byteaddress,
                                                std_2s60_burst_11_upstream_byteenable,
                                                std_2s60_burst_11_upstream_debugaccess,
                                                std_2s60_burst_11_upstream_read,
                                                std_2s60_burst_11_upstream_readdata_from_sa,
                                                std_2s60_burst_11_upstream_waitrequest_from_sa,
                                                std_2s60_burst_11_upstream_write,
                                                std_2s60_burst_11_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_11_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_11_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_11_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_11_upstream;
  output           d1_std_2s60_burst_11_upstream_end_xfer;
  output  [  2: 0] std_2s60_burst_11_upstream_address;
  output  [  3: 0] std_2s60_burst_11_upstream_burstcount;
  output  [  4: 0] std_2s60_burst_11_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_11_upstream_byteenable;
  output           std_2s60_burst_11_upstream_debugaccess;
  output           std_2s60_burst_11_upstream_read;
  output  [ 31: 0] std_2s60_burst_11_upstream_readdata_from_sa;
  output           std_2s60_burst_11_upstream_waitrequest_from_sa;
  output           std_2s60_burst_11_upstream_write;
  output  [ 31: 0] std_2s60_burst_11_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_11_upstream_readdata;
  input            std_2s60_burst_11_upstream_readdatavalid;
  input            std_2s60_burst_11_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_11_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_11_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_11_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_11_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_11_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_11_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_11_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_11_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_11_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_11_upstream_from_cpu_data_master;
  wire    [  2: 0] std_2s60_burst_11_upstream_address;
  wire             std_2s60_burst_11_upstream_allgrants;
  wire             std_2s60_burst_11_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_11_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_11_upstream_any_continuerequest;
  wire             std_2s60_burst_11_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_11_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_11_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_11_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_11_upstream_bbt_burstcounter;
  wire             std_2s60_burst_11_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_11_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_11_upstream_burstcount;
  wire             std_2s60_burst_11_upstream_burstcount_fifo_empty;
  wire    [  4: 0] std_2s60_burst_11_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_11_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_11_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_11_upstream_current_burst_minus_one;
  wire             std_2s60_burst_11_upstream_debugaccess;
  wire             std_2s60_burst_11_upstream_end_xfer;
  wire             std_2s60_burst_11_upstream_firsttransfer;
  wire             std_2s60_burst_11_upstream_grant_vector;
  wire             std_2s60_burst_11_upstream_in_a_read_cycle;
  wire             std_2s60_burst_11_upstream_in_a_write_cycle;
  reg              std_2s60_burst_11_upstream_load_fifo;
  wire             std_2s60_burst_11_upstream_master_qreq_vector;
  wire             std_2s60_burst_11_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_11_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_11_upstream_next_burst_count;
  wire             std_2s60_burst_11_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_11_upstream_read;
  wire    [ 31: 0] std_2s60_burst_11_upstream_readdata_from_sa;
  wire             std_2s60_burst_11_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_11_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_11_upstream_selected_burstcount;
  reg              std_2s60_burst_11_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_11_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_11_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_11_upstream_transaction_burst_count;
  wire             std_2s60_burst_11_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_11_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_11_upstream_waits_for_read;
  wire             std_2s60_burst_11_upstream_waits_for_write;
  wire             std_2s60_burst_11_upstream_write;
  wire    [ 31: 0] std_2s60_burst_11_upstream_writedata;
  wire             wait_for_std_2s60_burst_11_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_11_upstream_end_xfer;
    end


  assign std_2s60_burst_11_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_11_upstream));
  //assign std_2s60_burst_11_upstream_readdatavalid_from_sa = std_2s60_burst_11_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_11_upstream_readdatavalid_from_sa = std_2s60_burst_11_upstream_readdatavalid;

  //assign std_2s60_burst_11_upstream_readdata_from_sa = std_2s60_burst_11_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_11_upstream_readdata_from_sa = std_2s60_burst_11_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_11_upstream = ({cpu_data_master_address_to_slave[25 : 3] , 3'b0} == 26'h2131880) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_11_upstream_waitrequest_from_sa = std_2s60_burst_11_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_11_upstream_waitrequest_from_sa = std_2s60_burst_11_upstream_waitrequest;

  //std_2s60_burst_11_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_11_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_11_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_11_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_11_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_11_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_11_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_11_upstream;

  //std_2s60_burst_11_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_11_upstream_arb_share_counter_next_value = std_2s60_burst_11_upstream_firsttransfer ? (std_2s60_burst_11_upstream_arb_share_set_values - 1) : |std_2s60_burst_11_upstream_arb_share_counter ? (std_2s60_burst_11_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_11_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_11_upstream_allgrants = |std_2s60_burst_11_upstream_grant_vector;

  //std_2s60_burst_11_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_11_upstream_end_xfer = ~(std_2s60_burst_11_upstream_waits_for_read | std_2s60_burst_11_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream = std_2s60_burst_11_upstream_end_xfer & (~std_2s60_burst_11_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_11_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_11_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream & std_2s60_burst_11_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream & ~std_2s60_burst_11_upstream_non_bursting_master_requests);

  //std_2s60_burst_11_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_11_upstream_arb_counter_enable)
          std_2s60_burst_11_upstream_arb_share_counter <= std_2s60_burst_11_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_11_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_11_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_11_upstream & ~std_2s60_burst_11_upstream_non_bursting_master_requests))
          std_2s60_burst_11_upstream_slavearbiterlockenable <= |std_2s60_burst_11_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_11/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_11_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_11_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_11_upstream_slavearbiterlockenable2 = |std_2s60_burst_11_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_11/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_11_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_11_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_11_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_11_upstream = cpu_data_master_requests_std_2s60_burst_11_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_11_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_11_upstream_move_on_to_next_transaction = std_2s60_burst_11_upstream_this_cycle_is_the_last_burst & std_2s60_burst_11_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_11_upstream, which is an e_mux
  assign std_2s60_burst_11_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_11_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_11_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_11_upstream_module burstcount_fifo_for_std_2s60_burst_11_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_11_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_11_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_11_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_11_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read & std_2s60_burst_11_upstream_load_fifo & ~(std_2s60_burst_11_upstream_this_cycle_is_the_last_burst & std_2s60_burst_11_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_11_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_11_upstream_current_burst_minus_one = std_2s60_burst_11_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_11_upstream, which is an e_mux
  assign std_2s60_burst_11_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read) & ~std_2s60_burst_11_upstream_load_fifo))? std_2s60_burst_11_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read & std_2s60_burst_11_upstream_this_cycle_is_the_last_burst & std_2s60_burst_11_upstream_burstcount_fifo_empty))? std_2s60_burst_11_upstream_selected_burstcount :
    (std_2s60_burst_11_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_11_upstream_transaction_burst_count :
    std_2s60_burst_11_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_11_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_current_burst <= 0;
      else if (std_2s60_burst_11_upstream_readdatavalid_from_sa | (~std_2s60_burst_11_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read)))
          std_2s60_burst_11_upstream_current_burst <= std_2s60_burst_11_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_11_upstream_load_fifo = (~std_2s60_burst_11_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read) & std_2s60_burst_11_upstream_load_fifo))? 1 :
    ~std_2s60_burst_11_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read) & ~std_2s60_burst_11_upstream_load_fifo | std_2s60_burst_11_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_11_upstream_load_fifo <= p0_std_2s60_burst_11_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_11_upstream, which is an e_assign
  assign std_2s60_burst_11_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_11_upstream_current_burst_minus_one) & std_2s60_burst_11_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_11_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_11_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_11_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_11_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_11_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_11_upstream),
      .full                 (),
      .read                 (std_2s60_burst_11_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_11_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_11_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_11_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_11_upstream = std_2s60_burst_11_upstream_readdatavalid_from_sa;

  //std_2s60_burst_11_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_11_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_11/upstream, which is an e_mux
  assign std_2s60_burst_11_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_11_upstream = cpu_data_master_qualified_request_std_2s60_burst_11_upstream;

  //cpu/data_master saved-grant std_2s60_burst_11/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_11_upstream = cpu_data_master_requests_std_2s60_burst_11_upstream;

  //allow new arb cycle for std_2s60_burst_11/upstream, which is an e_assign
  assign std_2s60_burst_11_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_11_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_11_upstream_master_qreq_vector = 1;

  //std_2s60_burst_11_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_11_upstream_firsttransfer = std_2s60_burst_11_upstream_begins_xfer ? std_2s60_burst_11_upstream_unreg_firsttransfer : std_2s60_burst_11_upstream_reg_firsttransfer;

  //std_2s60_burst_11_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_11_upstream_unreg_firsttransfer = ~(std_2s60_burst_11_upstream_slavearbiterlockenable & std_2s60_burst_11_upstream_any_continuerequest);

  //std_2s60_burst_11_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_11_upstream_begins_xfer)
          std_2s60_burst_11_upstream_reg_firsttransfer <= std_2s60_burst_11_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_11_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_11_upstream_next_bbt_burstcount = ((((std_2s60_burst_11_upstream_write) && (std_2s60_burst_11_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_11_upstream_burstcount - 1) :
    ((((std_2s60_burst_11_upstream_read) && (std_2s60_burst_11_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_11_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_11_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_11_upstream_begins_xfer)
          std_2s60_burst_11_upstream_bbt_burstcounter <= std_2s60_burst_11_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_11_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_11_upstream_beginbursttransfer_internal = std_2s60_burst_11_upstream_begins_xfer & (std_2s60_burst_11_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_11_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_11_upstream_read = cpu_data_master_granted_std_2s60_burst_11_upstream & cpu_data_master_read;

  //std_2s60_burst_11_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_11_upstream_write = cpu_data_master_granted_std_2s60_burst_11_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_11_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_11_upstream_address mux, which is an e_mux
  assign std_2s60_burst_11_upstream_address = shifted_address_to_std_2s60_burst_11_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_11_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_11_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_11_upstream_end_xfer <= std_2s60_burst_11_upstream_end_xfer;
    end


  //std_2s60_burst_11_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_11_upstream_waits_for_read = std_2s60_burst_11_upstream_in_a_read_cycle & std_2s60_burst_11_upstream_waitrequest_from_sa;

  //std_2s60_burst_11_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_11_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_11_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_11_upstream_in_a_read_cycle;

  //std_2s60_burst_11_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_11_upstream_waits_for_write = std_2s60_burst_11_upstream_in_a_write_cycle & std_2s60_burst_11_upstream_waitrequest_from_sa;

  //std_2s60_burst_11_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_11_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_11_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_11_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_11_upstream_counter = 0;
  //std_2s60_burst_11_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_11_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_11_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_11_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_11_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_11_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_11_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_11/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_11_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_11/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_11_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                  jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                  jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                  reset_n,
                                                  std_2s60_burst_11_downstream_address,
                                                  std_2s60_burst_11_downstream_burstcount,
                                                  std_2s60_burst_11_downstream_byteenable,
                                                  std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave,
                                                  std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave,
                                                  std_2s60_burst_11_downstream_read,
                                                  std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                  std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave,
                                                  std_2s60_burst_11_downstream_write,
                                                  std_2s60_burst_11_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_11_downstream_address_to_slave,
                                                  std_2s60_burst_11_downstream_latency_counter,
                                                  std_2s60_burst_11_downstream_readdata,
                                                  std_2s60_burst_11_downstream_readdatavalid,
                                                  std_2s60_burst_11_downstream_reset_n,
                                                  std_2s60_burst_11_downstream_waitrequest
                                               )
;

  output  [  2: 0] std_2s60_burst_11_downstream_address_to_slave;
  output           std_2s60_burst_11_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_11_downstream_readdata;
  output           std_2s60_burst_11_downstream_readdatavalid;
  output           std_2s60_burst_11_downstream_reset_n;
  output           std_2s60_burst_11_downstream_waitrequest;
  input            clk;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input            reset_n;
  input   [  2: 0] std_2s60_burst_11_downstream_address;
  input            std_2s60_burst_11_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_11_downstream_byteenable;
  input            std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave;
  input            std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  input            std_2s60_burst_11_downstream_read;
  input            std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave;
  input            std_2s60_burst_11_downstream_write;
  input   [ 31: 0] std_2s60_burst_11_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             pre_flush_std_2s60_burst_11_downstream_readdatavalid;
  wire             r_0;
  reg     [  2: 0] std_2s60_burst_11_downstream_address_last_time;
  wire    [  2: 0] std_2s60_burst_11_downstream_address_to_slave;
  reg              std_2s60_burst_11_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_11_downstream_byteenable_last_time;
  wire             std_2s60_burst_11_downstream_latency_counter;
  reg              std_2s60_burst_11_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_11_downstream_readdata;
  wire             std_2s60_burst_11_downstream_readdatavalid;
  wire             std_2s60_burst_11_downstream_reset_n;
  wire             std_2s60_burst_11_downstream_run;
  wire             std_2s60_burst_11_downstream_waitrequest;
  reg              std_2s60_burst_11_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_11_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave | ~std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave) & ((~std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave | ~(std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write)))) & ((~std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave | ~(std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_11_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_11_downstream_address_to_slave = std_2s60_burst_11_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_11_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_11_downstream_readdatavalid = 0 |
    pre_flush_std_2s60_burst_11_downstream_readdatavalid |
    std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave;

  //std_2s60_burst_11/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_11_downstream_readdata = jtag_uart_avalon_jtag_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_11_downstream_waitrequest = ~std_2s60_burst_11_downstream_run;

  //latent max counter, which is an e_assign
  assign std_2s60_burst_11_downstream_latency_counter = 0;

  //std_2s60_burst_11_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_11_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_11_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_address_last_time <= std_2s60_burst_11_downstream_address;
    end


  //std_2s60_burst_11/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_11_downstream_waitrequest & (std_2s60_burst_11_downstream_read | std_2s60_burst_11_downstream_write);
    end


  //std_2s60_burst_11_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_address != std_2s60_burst_11_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_11_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_burstcount_last_time <= std_2s60_burst_11_downstream_burstcount;
    end


  //std_2s60_burst_11_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_burstcount != std_2s60_burst_11_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_11_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_byteenable_last_time <= std_2s60_burst_11_downstream_byteenable;
    end


  //std_2s60_burst_11_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_byteenable != std_2s60_burst_11_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_11_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_read_last_time <= std_2s60_burst_11_downstream_read;
    end


  //std_2s60_burst_11_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_read != std_2s60_burst_11_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_11_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_write_last_time <= std_2s60_burst_11_downstream_write;
    end


  //std_2s60_burst_11_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_write != std_2s60_burst_11_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_11_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_11_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_11_downstream_writedata_last_time <= std_2s60_burst_11_downstream_writedata;
    end


  //std_2s60_burst_11_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_11_downstream_writedata != std_2s60_burst_11_downstream_writedata_last_time) & std_2s60_burst_11_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_11_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_12_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_12_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_12_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_12_upstream_readdata,
                                                std_2s60_burst_12_upstream_readdatavalid,
                                                std_2s60_burst_12_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_12_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_12_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_12_upstream,
                                                d1_std_2s60_burst_12_upstream_end_xfer,
                                                std_2s60_burst_12_upstream_address,
                                                std_2s60_burst_12_upstream_burstcount,
                                                std_2s60_burst_12_upstream_byteaddress,
                                                std_2s60_burst_12_upstream_byteenable,
                                                std_2s60_burst_12_upstream_debugaccess,
                                                std_2s60_burst_12_upstream_read,
                                                std_2s60_burst_12_upstream_readdata_from_sa,
                                                std_2s60_burst_12_upstream_waitrequest_from_sa,
                                                std_2s60_burst_12_upstream_write,
                                                std_2s60_burst_12_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_12_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_12_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_12_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_12_upstream;
  output           d1_std_2s60_burst_12_upstream_end_xfer;
  output  [  3: 0] std_2s60_burst_12_upstream_address;
  output  [  3: 0] std_2s60_burst_12_upstream_burstcount;
  output  [  4: 0] std_2s60_burst_12_upstream_byteaddress;
  output  [  1: 0] std_2s60_burst_12_upstream_byteenable;
  output           std_2s60_burst_12_upstream_debugaccess;
  output           std_2s60_burst_12_upstream_read;
  output  [ 15: 0] std_2s60_burst_12_upstream_readdata_from_sa;
  output           std_2s60_burst_12_upstream_waitrequest_from_sa;
  output           std_2s60_burst_12_upstream_write;
  output  [ 15: 0] std_2s60_burst_12_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_12_upstream_readdata;
  input            std_2s60_burst_12_upstream_readdatavalid;
  input            std_2s60_burst_12_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_12_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_12_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_12_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_12_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_12_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_12_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_12_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_12_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_12_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_12_upstream_from_cpu_data_master;
  wire    [  3: 0] std_2s60_burst_12_upstream_address;
  wire             std_2s60_burst_12_upstream_allgrants;
  wire             std_2s60_burst_12_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_12_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_12_upstream_any_continuerequest;
  wire             std_2s60_burst_12_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_12_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_12_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_12_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_12_upstream_bbt_burstcounter;
  wire             std_2s60_burst_12_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_12_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_12_upstream_burstcount;
  wire             std_2s60_burst_12_upstream_burstcount_fifo_empty;
  wire    [  4: 0] std_2s60_burst_12_upstream_byteaddress;
  wire    [  1: 0] std_2s60_burst_12_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_12_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_12_upstream_current_burst_minus_one;
  wire             std_2s60_burst_12_upstream_debugaccess;
  wire             std_2s60_burst_12_upstream_end_xfer;
  wire             std_2s60_burst_12_upstream_firsttransfer;
  wire             std_2s60_burst_12_upstream_grant_vector;
  wire             std_2s60_burst_12_upstream_in_a_read_cycle;
  wire             std_2s60_burst_12_upstream_in_a_write_cycle;
  reg              std_2s60_burst_12_upstream_load_fifo;
  wire             std_2s60_burst_12_upstream_master_qreq_vector;
  wire             std_2s60_burst_12_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_12_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_12_upstream_next_burst_count;
  wire             std_2s60_burst_12_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_12_upstream_read;
  wire    [ 15: 0] std_2s60_burst_12_upstream_readdata_from_sa;
  wire             std_2s60_burst_12_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_12_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_12_upstream_selected_burstcount;
  reg              std_2s60_burst_12_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_12_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_12_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_12_upstream_transaction_burst_count;
  wire             std_2s60_burst_12_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_12_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_12_upstream_waits_for_read;
  wire             std_2s60_burst_12_upstream_waits_for_write;
  wire             std_2s60_burst_12_upstream_write;
  wire    [ 15: 0] std_2s60_burst_12_upstream_writedata;
  wire             wait_for_std_2s60_burst_12_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_12_upstream_end_xfer;
    end


  assign std_2s60_burst_12_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_12_upstream));
  //assign std_2s60_burst_12_upstream_readdatavalid_from_sa = std_2s60_burst_12_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_12_upstream_readdatavalid_from_sa = std_2s60_burst_12_upstream_readdatavalid;

  //assign std_2s60_burst_12_upstream_readdata_from_sa = std_2s60_burst_12_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_12_upstream_readdata_from_sa = std_2s60_burst_12_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_12_upstream = ({cpu_data_master_address_to_slave[25 : 5] , 5'b0} == 26'h2131820) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_12_upstream_waitrequest_from_sa = std_2s60_burst_12_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_12_upstream_waitrequest_from_sa = std_2s60_burst_12_upstream_waitrequest;

  //std_2s60_burst_12_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_12_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_12_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_12_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_12_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_12_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_12_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_12_upstream;

  //std_2s60_burst_12_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_12_upstream_arb_share_counter_next_value = std_2s60_burst_12_upstream_firsttransfer ? (std_2s60_burst_12_upstream_arb_share_set_values - 1) : |std_2s60_burst_12_upstream_arb_share_counter ? (std_2s60_burst_12_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_12_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_12_upstream_allgrants = |std_2s60_burst_12_upstream_grant_vector;

  //std_2s60_burst_12_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_12_upstream_end_xfer = ~(std_2s60_burst_12_upstream_waits_for_read | std_2s60_burst_12_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream = std_2s60_burst_12_upstream_end_xfer & (~std_2s60_burst_12_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_12_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_12_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream & std_2s60_burst_12_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream & ~std_2s60_burst_12_upstream_non_bursting_master_requests);

  //std_2s60_burst_12_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_12_upstream_arb_counter_enable)
          std_2s60_burst_12_upstream_arb_share_counter <= std_2s60_burst_12_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_12_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_12_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_12_upstream & ~std_2s60_burst_12_upstream_non_bursting_master_requests))
          std_2s60_burst_12_upstream_slavearbiterlockenable <= |std_2s60_burst_12_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_12/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_12_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_12_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_12_upstream_slavearbiterlockenable2 = |std_2s60_burst_12_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_12/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_12_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_12_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_12_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_12_upstream = cpu_data_master_requests_std_2s60_burst_12_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_12_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_12_upstream_move_on_to_next_transaction = std_2s60_burst_12_upstream_this_cycle_is_the_last_burst & std_2s60_burst_12_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_12_upstream, which is an e_mux
  assign std_2s60_burst_12_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_12_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_12_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_12_upstream_module burstcount_fifo_for_std_2s60_burst_12_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_12_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_12_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_12_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_12_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read & std_2s60_burst_12_upstream_load_fifo & ~(std_2s60_burst_12_upstream_this_cycle_is_the_last_burst & std_2s60_burst_12_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_12_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_12_upstream_current_burst_minus_one = std_2s60_burst_12_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_12_upstream, which is an e_mux
  assign std_2s60_burst_12_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read) & ~std_2s60_burst_12_upstream_load_fifo))? std_2s60_burst_12_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read & std_2s60_burst_12_upstream_this_cycle_is_the_last_burst & std_2s60_burst_12_upstream_burstcount_fifo_empty))? std_2s60_burst_12_upstream_selected_burstcount :
    (std_2s60_burst_12_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_12_upstream_transaction_burst_count :
    std_2s60_burst_12_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_12_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_current_burst <= 0;
      else if (std_2s60_burst_12_upstream_readdatavalid_from_sa | (~std_2s60_burst_12_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read)))
          std_2s60_burst_12_upstream_current_burst <= std_2s60_burst_12_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_12_upstream_load_fifo = (~std_2s60_burst_12_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read) & std_2s60_burst_12_upstream_load_fifo))? 1 :
    ~std_2s60_burst_12_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read) & ~std_2s60_burst_12_upstream_load_fifo | std_2s60_burst_12_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_12_upstream_load_fifo <= p0_std_2s60_burst_12_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_12_upstream, which is an e_assign
  assign std_2s60_burst_12_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_12_upstream_current_burst_minus_one) & std_2s60_burst_12_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_12_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_12_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_12_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_12_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_12_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_12_upstream),
      .full                 (),
      .read                 (std_2s60_burst_12_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_12_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_12_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_12_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_12_upstream = std_2s60_burst_12_upstream_readdatavalid_from_sa;

  //std_2s60_burst_12_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_12_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_12/upstream, which is an e_mux
  assign std_2s60_burst_12_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_12_upstream = cpu_data_master_qualified_request_std_2s60_burst_12_upstream;

  //cpu/data_master saved-grant std_2s60_burst_12/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_12_upstream = cpu_data_master_requests_std_2s60_burst_12_upstream;

  //allow new arb cycle for std_2s60_burst_12/upstream, which is an e_assign
  assign std_2s60_burst_12_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_12_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_12_upstream_master_qreq_vector = 1;

  //std_2s60_burst_12_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_12_upstream_firsttransfer = std_2s60_burst_12_upstream_begins_xfer ? std_2s60_burst_12_upstream_unreg_firsttransfer : std_2s60_burst_12_upstream_reg_firsttransfer;

  //std_2s60_burst_12_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_12_upstream_unreg_firsttransfer = ~(std_2s60_burst_12_upstream_slavearbiterlockenable & std_2s60_burst_12_upstream_any_continuerequest);

  //std_2s60_burst_12_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_12_upstream_begins_xfer)
          std_2s60_burst_12_upstream_reg_firsttransfer <= std_2s60_burst_12_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_12_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_12_upstream_next_bbt_burstcount = ((((std_2s60_burst_12_upstream_write) && (std_2s60_burst_12_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_12_upstream_burstcount - 1) :
    ((((std_2s60_burst_12_upstream_read) && (std_2s60_burst_12_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_12_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_12_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_12_upstream_begins_xfer)
          std_2s60_burst_12_upstream_bbt_burstcounter <= std_2s60_burst_12_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_12_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_12_upstream_beginbursttransfer_internal = std_2s60_burst_12_upstream_begins_xfer & (std_2s60_burst_12_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_12_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_12_upstream_read = cpu_data_master_granted_std_2s60_burst_12_upstream & cpu_data_master_read;

  //std_2s60_burst_12_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_12_upstream_write = cpu_data_master_granted_std_2s60_burst_12_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_12_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_12_upstream_address mux, which is an e_mux
  assign std_2s60_burst_12_upstream_address = shifted_address_to_std_2s60_burst_12_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_12_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_12_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_12_upstream_end_xfer <= std_2s60_burst_12_upstream_end_xfer;
    end


  //std_2s60_burst_12_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_12_upstream_waits_for_read = std_2s60_burst_12_upstream_in_a_read_cycle & std_2s60_burst_12_upstream_waitrequest_from_sa;

  //std_2s60_burst_12_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_12_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_12_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_12_upstream_in_a_read_cycle;

  //std_2s60_burst_12_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_12_upstream_waits_for_write = std_2s60_burst_12_upstream_in_a_write_cycle & std_2s60_burst_12_upstream_waitrequest_from_sa;

  //std_2s60_burst_12_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_12_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_12_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_12_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_12_upstream_counter = 0;
  //std_2s60_burst_12_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_12_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_12_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_12_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_12_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_12_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_12_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_12/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_12_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_12/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_12_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_high_res_timer_s1_end_xfer,
                                                  high_res_timer_s1_readdata_from_sa,
                                                  reset_n,
                                                  std_2s60_burst_12_downstream_address,
                                                  std_2s60_burst_12_downstream_burstcount,
                                                  std_2s60_burst_12_downstream_byteenable,
                                                  std_2s60_burst_12_downstream_granted_high_res_timer_s1,
                                                  std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1,
                                                  std_2s60_burst_12_downstream_read,
                                                  std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1,
                                                  std_2s60_burst_12_downstream_requests_high_res_timer_s1,
                                                  std_2s60_burst_12_downstream_write,
                                                  std_2s60_burst_12_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_12_downstream_address_to_slave,
                                                  std_2s60_burst_12_downstream_latency_counter,
                                                  std_2s60_burst_12_downstream_readdata,
                                                  std_2s60_burst_12_downstream_readdatavalid,
                                                  std_2s60_burst_12_downstream_reset_n,
                                                  std_2s60_burst_12_downstream_waitrequest
                                               )
;

  output  [  3: 0] std_2s60_burst_12_downstream_address_to_slave;
  output           std_2s60_burst_12_downstream_latency_counter;
  output  [ 15: 0] std_2s60_burst_12_downstream_readdata;
  output           std_2s60_burst_12_downstream_readdatavalid;
  output           std_2s60_burst_12_downstream_reset_n;
  output           std_2s60_burst_12_downstream_waitrequest;
  input            clk;
  input            d1_high_res_timer_s1_end_xfer;
  input   [ 15: 0] high_res_timer_s1_readdata_from_sa;
  input            reset_n;
  input   [  3: 0] std_2s60_burst_12_downstream_address;
  input            std_2s60_burst_12_downstream_burstcount;
  input   [  1: 0] std_2s60_burst_12_downstream_byteenable;
  input            std_2s60_burst_12_downstream_granted_high_res_timer_s1;
  input            std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1;
  input            std_2s60_burst_12_downstream_read;
  input            std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1;
  input            std_2s60_burst_12_downstream_requests_high_res_timer_s1;
  input            std_2s60_burst_12_downstream_write;
  input   [ 15: 0] std_2s60_burst_12_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             pre_flush_std_2s60_burst_12_downstream_readdatavalid;
  wire             r_0;
  reg     [  3: 0] std_2s60_burst_12_downstream_address_last_time;
  wire    [  3: 0] std_2s60_burst_12_downstream_address_to_slave;
  reg              std_2s60_burst_12_downstream_burstcount_last_time;
  reg     [  1: 0] std_2s60_burst_12_downstream_byteenable_last_time;
  wire             std_2s60_burst_12_downstream_latency_counter;
  reg              std_2s60_burst_12_downstream_read_last_time;
  wire    [ 15: 0] std_2s60_burst_12_downstream_readdata;
  wire             std_2s60_burst_12_downstream_readdatavalid;
  wire             std_2s60_burst_12_downstream_reset_n;
  wire             std_2s60_burst_12_downstream_run;
  wire             std_2s60_burst_12_downstream_waitrequest;
  reg              std_2s60_burst_12_downstream_write_last_time;
  reg     [ 15: 0] std_2s60_burst_12_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 | ~std_2s60_burst_12_downstream_requests_high_res_timer_s1) & ((~std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 | ~std_2s60_burst_12_downstream_read | (1 & ~d1_high_res_timer_s1_end_xfer & std_2s60_burst_12_downstream_read))) & ((~std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 | ~std_2s60_burst_12_downstream_write | (1 & std_2s60_burst_12_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_12_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_12_downstream_address_to_slave = std_2s60_burst_12_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_12_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_12_downstream_readdatavalid = 0 |
    pre_flush_std_2s60_burst_12_downstream_readdatavalid |
    std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1;

  //std_2s60_burst_12/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_12_downstream_readdata = high_res_timer_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_12_downstream_waitrequest = ~std_2s60_burst_12_downstream_run;

  //latent max counter, which is an e_assign
  assign std_2s60_burst_12_downstream_latency_counter = 0;

  //std_2s60_burst_12_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_12_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_12_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_address_last_time <= std_2s60_burst_12_downstream_address;
    end


  //std_2s60_burst_12/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_12_downstream_waitrequest & (std_2s60_burst_12_downstream_read | std_2s60_burst_12_downstream_write);
    end


  //std_2s60_burst_12_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_address != std_2s60_burst_12_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_12_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_burstcount_last_time <= std_2s60_burst_12_downstream_burstcount;
    end


  //std_2s60_burst_12_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_burstcount != std_2s60_burst_12_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_12_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_byteenable_last_time <= std_2s60_burst_12_downstream_byteenable;
    end


  //std_2s60_burst_12_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_byteenable != std_2s60_burst_12_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_12_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_read_last_time <= std_2s60_burst_12_downstream_read;
    end


  //std_2s60_burst_12_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_read != std_2s60_burst_12_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_12_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_write_last_time <= std_2s60_burst_12_downstream_write;
    end


  //std_2s60_burst_12_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_write != std_2s60_burst_12_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_12_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_12_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_12_downstream_writedata_last_time <= std_2s60_burst_12_downstream_writedata;
    end


  //std_2s60_burst_12_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_12_downstream_writedata != std_2s60_burst_12_downstream_writedata_last_time) & std_2s60_burst_12_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_12_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_13_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_13_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_13_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_13_upstream_readdata,
                                                std_2s60_burst_13_upstream_readdatavalid,
                                                std_2s60_burst_13_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_13_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_13_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_13_upstream,
                                                d1_std_2s60_burst_13_upstream_end_xfer,
                                                std_2s60_burst_13_upstream_address,
                                                std_2s60_burst_13_upstream_burstcount,
                                                std_2s60_burst_13_upstream_byteaddress,
                                                std_2s60_burst_13_upstream_byteenable,
                                                std_2s60_burst_13_upstream_debugaccess,
                                                std_2s60_burst_13_upstream_read,
                                                std_2s60_burst_13_upstream_readdata_from_sa,
                                                std_2s60_burst_13_upstream_waitrequest_from_sa,
                                                std_2s60_burst_13_upstream_write,
                                                std_2s60_burst_13_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_13_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_13_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_13_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_13_upstream;
  output           d1_std_2s60_burst_13_upstream_end_xfer;
  output  [  1: 0] std_2s60_burst_13_upstream_address;
  output  [  3: 0] std_2s60_burst_13_upstream_burstcount;
  output  [  1: 0] std_2s60_burst_13_upstream_byteaddress;
  output           std_2s60_burst_13_upstream_byteenable;
  output           std_2s60_burst_13_upstream_debugaccess;
  output           std_2s60_burst_13_upstream_read;
  output  [  7: 0] std_2s60_burst_13_upstream_readdata_from_sa;
  output           std_2s60_burst_13_upstream_waitrequest_from_sa;
  output           std_2s60_burst_13_upstream_write;
  output  [  7: 0] std_2s60_burst_13_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [  7: 0] std_2s60_burst_13_upstream_readdata;
  input            std_2s60_burst_13_upstream_readdatavalid;
  input            std_2s60_burst_13_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_13_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_13_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_13_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_13_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_13_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_13_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_13_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_13_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_13_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_13_upstream_from_cpu_data_master;
  wire    [  1: 0] std_2s60_burst_13_upstream_address;
  wire             std_2s60_burst_13_upstream_allgrants;
  wire             std_2s60_burst_13_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_13_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_13_upstream_any_continuerequest;
  wire             std_2s60_burst_13_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_13_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_13_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_13_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_13_upstream_bbt_burstcounter;
  wire             std_2s60_burst_13_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_13_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_13_upstream_burstcount;
  wire             std_2s60_burst_13_upstream_burstcount_fifo_empty;
  wire    [  1: 0] std_2s60_burst_13_upstream_byteaddress;
  wire             std_2s60_burst_13_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_13_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_13_upstream_current_burst_minus_one;
  wire             std_2s60_burst_13_upstream_debugaccess;
  wire             std_2s60_burst_13_upstream_end_xfer;
  wire             std_2s60_burst_13_upstream_firsttransfer;
  wire             std_2s60_burst_13_upstream_grant_vector;
  wire             std_2s60_burst_13_upstream_in_a_read_cycle;
  wire             std_2s60_burst_13_upstream_in_a_write_cycle;
  reg              std_2s60_burst_13_upstream_load_fifo;
  wire             std_2s60_burst_13_upstream_master_qreq_vector;
  wire             std_2s60_burst_13_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_13_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_13_upstream_next_burst_count;
  wire             std_2s60_burst_13_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_13_upstream_read;
  wire    [  7: 0] std_2s60_burst_13_upstream_readdata_from_sa;
  wire             std_2s60_burst_13_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_13_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_13_upstream_selected_burstcount;
  reg              std_2s60_burst_13_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_13_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_13_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_13_upstream_transaction_burst_count;
  wire             std_2s60_burst_13_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_13_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_13_upstream_waits_for_read;
  wire             std_2s60_burst_13_upstream_waits_for_write;
  wire             std_2s60_burst_13_upstream_write;
  wire    [  7: 0] std_2s60_burst_13_upstream_writedata;
  wire             wait_for_std_2s60_burst_13_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_13_upstream_end_xfer;
    end


  assign std_2s60_burst_13_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_13_upstream));
  //assign std_2s60_burst_13_upstream_readdatavalid_from_sa = std_2s60_burst_13_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_13_upstream_readdatavalid_from_sa = std_2s60_burst_13_upstream_readdatavalid;

  //assign std_2s60_burst_13_upstream_readdata_from_sa = std_2s60_burst_13_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_13_upstream_readdata_from_sa = std_2s60_burst_13_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_13_upstream = ({cpu_data_master_address_to_slave[25 : 4] , 4'b0} == 26'h2131870) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_13_upstream_waitrequest_from_sa = std_2s60_burst_13_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_13_upstream_waitrequest_from_sa = std_2s60_burst_13_upstream_waitrequest;

  //std_2s60_burst_13_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_13_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_13_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_13_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_13_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_13_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_13_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_13_upstream;

  //std_2s60_burst_13_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_13_upstream_arb_share_counter_next_value = std_2s60_burst_13_upstream_firsttransfer ? (std_2s60_burst_13_upstream_arb_share_set_values - 1) : |std_2s60_burst_13_upstream_arb_share_counter ? (std_2s60_burst_13_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_13_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_13_upstream_allgrants = |std_2s60_burst_13_upstream_grant_vector;

  //std_2s60_burst_13_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_13_upstream_end_xfer = ~(std_2s60_burst_13_upstream_waits_for_read | std_2s60_burst_13_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream = std_2s60_burst_13_upstream_end_xfer & (~std_2s60_burst_13_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_13_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_13_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream & std_2s60_burst_13_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream & ~std_2s60_burst_13_upstream_non_bursting_master_requests);

  //std_2s60_burst_13_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_13_upstream_arb_counter_enable)
          std_2s60_burst_13_upstream_arb_share_counter <= std_2s60_burst_13_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_13_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_13_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_13_upstream & ~std_2s60_burst_13_upstream_non_bursting_master_requests))
          std_2s60_burst_13_upstream_slavearbiterlockenable <= |std_2s60_burst_13_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_13/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_13_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_13_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_13_upstream_slavearbiterlockenable2 = |std_2s60_burst_13_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_13/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_13_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_13_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_13_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_13_upstream = cpu_data_master_requests_std_2s60_burst_13_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_13_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_13_upstream_move_on_to_next_transaction = std_2s60_burst_13_upstream_this_cycle_is_the_last_burst & std_2s60_burst_13_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_13_upstream, which is an e_mux
  assign std_2s60_burst_13_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_13_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_13_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_13_upstream_module burstcount_fifo_for_std_2s60_burst_13_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_13_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_13_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_13_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_13_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read & std_2s60_burst_13_upstream_load_fifo & ~(std_2s60_burst_13_upstream_this_cycle_is_the_last_burst & std_2s60_burst_13_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_13_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_13_upstream_current_burst_minus_one = std_2s60_burst_13_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_13_upstream, which is an e_mux
  assign std_2s60_burst_13_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read) & ~std_2s60_burst_13_upstream_load_fifo))? std_2s60_burst_13_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read & std_2s60_burst_13_upstream_this_cycle_is_the_last_burst & std_2s60_burst_13_upstream_burstcount_fifo_empty))? std_2s60_burst_13_upstream_selected_burstcount :
    (std_2s60_burst_13_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_13_upstream_transaction_burst_count :
    std_2s60_burst_13_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_13_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_current_burst <= 0;
      else if (std_2s60_burst_13_upstream_readdatavalid_from_sa | (~std_2s60_burst_13_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read)))
          std_2s60_burst_13_upstream_current_burst <= std_2s60_burst_13_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_13_upstream_load_fifo = (~std_2s60_burst_13_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read) & std_2s60_burst_13_upstream_load_fifo))? 1 :
    ~std_2s60_burst_13_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read) & ~std_2s60_burst_13_upstream_load_fifo | std_2s60_burst_13_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_13_upstream_load_fifo <= p0_std_2s60_burst_13_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_13_upstream, which is an e_assign
  assign std_2s60_burst_13_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_13_upstream_current_burst_minus_one) & std_2s60_burst_13_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_13_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_13_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_13_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_13_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_13_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_13_upstream),
      .full                 (),
      .read                 (std_2s60_burst_13_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_13_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_13_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_13_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_13_upstream = std_2s60_burst_13_upstream_readdatavalid_from_sa;

  //std_2s60_burst_13_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_13_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_13/upstream, which is an e_mux
  assign std_2s60_burst_13_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_13_upstream = cpu_data_master_qualified_request_std_2s60_burst_13_upstream;

  //cpu/data_master saved-grant std_2s60_burst_13/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_13_upstream = cpu_data_master_requests_std_2s60_burst_13_upstream;

  //allow new arb cycle for std_2s60_burst_13/upstream, which is an e_assign
  assign std_2s60_burst_13_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_13_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_13_upstream_master_qreq_vector = 1;

  //std_2s60_burst_13_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_13_upstream_firsttransfer = std_2s60_burst_13_upstream_begins_xfer ? std_2s60_burst_13_upstream_unreg_firsttransfer : std_2s60_burst_13_upstream_reg_firsttransfer;

  //std_2s60_burst_13_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_13_upstream_unreg_firsttransfer = ~(std_2s60_burst_13_upstream_slavearbiterlockenable & std_2s60_burst_13_upstream_any_continuerequest);

  //std_2s60_burst_13_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_13_upstream_begins_xfer)
          std_2s60_burst_13_upstream_reg_firsttransfer <= std_2s60_burst_13_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_13_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_13_upstream_next_bbt_burstcount = ((((std_2s60_burst_13_upstream_write) && (std_2s60_burst_13_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_13_upstream_burstcount - 1) :
    ((((std_2s60_burst_13_upstream_read) && (std_2s60_burst_13_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_13_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_13_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_13_upstream_begins_xfer)
          std_2s60_burst_13_upstream_bbt_burstcounter <= std_2s60_burst_13_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_13_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_13_upstream_beginbursttransfer_internal = std_2s60_burst_13_upstream_begins_xfer & (std_2s60_burst_13_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_13_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_13_upstream_read = cpu_data_master_granted_std_2s60_burst_13_upstream & cpu_data_master_read;

  //std_2s60_burst_13_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_13_upstream_write = cpu_data_master_granted_std_2s60_burst_13_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_13_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_13_upstream_address mux, which is an e_mux
  assign std_2s60_burst_13_upstream_address = shifted_address_to_std_2s60_burst_13_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_13_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_13_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_13_upstream_end_xfer <= std_2s60_burst_13_upstream_end_xfer;
    end


  //std_2s60_burst_13_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_13_upstream_waits_for_read = std_2s60_burst_13_upstream_in_a_read_cycle & std_2s60_burst_13_upstream_waitrequest_from_sa;

  //std_2s60_burst_13_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_13_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_13_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_13_upstream_in_a_read_cycle;

  //std_2s60_burst_13_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_13_upstream_waits_for_write = std_2s60_burst_13_upstream_in_a_write_cycle & std_2s60_burst_13_upstream_waitrequest_from_sa;

  //std_2s60_burst_13_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_13_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_13_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_13_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_13_upstream_counter = 0;
  //std_2s60_burst_13_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_13_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_13_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_13_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_13_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_13_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_13_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_13/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_13_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_13/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_13_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_reconfig_request_pio_s1_end_xfer,
                                                  reconfig_request_pio_s1_readdata_from_sa,
                                                  reset_n,
                                                  std_2s60_burst_13_downstream_address,
                                                  std_2s60_burst_13_downstream_burstcount,
                                                  std_2s60_burst_13_downstream_byteenable,
                                                  std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1,
                                                  std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1,
                                                  std_2s60_burst_13_downstream_read,
                                                  std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1,
                                                  std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1,
                                                  std_2s60_burst_13_downstream_write,
                                                  std_2s60_burst_13_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_13_downstream_address_to_slave,
                                                  std_2s60_burst_13_downstream_latency_counter,
                                                  std_2s60_burst_13_downstream_readdata,
                                                  std_2s60_burst_13_downstream_readdatavalid,
                                                  std_2s60_burst_13_downstream_reset_n,
                                                  std_2s60_burst_13_downstream_waitrequest
                                               )
;

  output  [  1: 0] std_2s60_burst_13_downstream_address_to_slave;
  output           std_2s60_burst_13_downstream_latency_counter;
  output  [  7: 0] std_2s60_burst_13_downstream_readdata;
  output           std_2s60_burst_13_downstream_readdatavalid;
  output           std_2s60_burst_13_downstream_reset_n;
  output           std_2s60_burst_13_downstream_waitrequest;
  input            clk;
  input            d1_reconfig_request_pio_s1_end_xfer;
  input            reconfig_request_pio_s1_readdata_from_sa;
  input            reset_n;
  input   [  1: 0] std_2s60_burst_13_downstream_address;
  input            std_2s60_burst_13_downstream_burstcount;
  input            std_2s60_burst_13_downstream_byteenable;
  input            std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1;
  input            std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1;
  input            std_2s60_burst_13_downstream_read;
  input            std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1;
  input            std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1;
  input            std_2s60_burst_13_downstream_write;
  input   [  7: 0] std_2s60_burst_13_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             pre_flush_std_2s60_burst_13_downstream_readdatavalid;
  wire             r_0;
  reg     [  1: 0] std_2s60_burst_13_downstream_address_last_time;
  wire    [  1: 0] std_2s60_burst_13_downstream_address_to_slave;
  reg              std_2s60_burst_13_downstream_burstcount_last_time;
  reg              std_2s60_burst_13_downstream_byteenable_last_time;
  wire             std_2s60_burst_13_downstream_latency_counter;
  reg              std_2s60_burst_13_downstream_read_last_time;
  wire    [  7: 0] std_2s60_burst_13_downstream_readdata;
  wire             std_2s60_burst_13_downstream_readdatavalid;
  wire             std_2s60_burst_13_downstream_reset_n;
  wire             std_2s60_burst_13_downstream_run;
  wire             std_2s60_burst_13_downstream_waitrequest;
  reg              std_2s60_burst_13_downstream_write_last_time;
  reg     [  7: 0] std_2s60_burst_13_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 | ~std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1) & ((~std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 | ~std_2s60_burst_13_downstream_read | (1 & ~d1_reconfig_request_pio_s1_end_xfer & std_2s60_burst_13_downstream_read))) & ((~std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 | ~std_2s60_burst_13_downstream_write | (1 & std_2s60_burst_13_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_13_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_13_downstream_address_to_slave = std_2s60_burst_13_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_13_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_13_downstream_readdatavalid = 0 |
    pre_flush_std_2s60_burst_13_downstream_readdatavalid |
    std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1;

  //std_2s60_burst_13/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_13_downstream_readdata = reconfig_request_pio_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_13_downstream_waitrequest = ~std_2s60_burst_13_downstream_run;

  //latent max counter, which is an e_assign
  assign std_2s60_burst_13_downstream_latency_counter = 0;

  //std_2s60_burst_13_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_13_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_13_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_address_last_time <= std_2s60_burst_13_downstream_address;
    end


  //std_2s60_burst_13/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_13_downstream_waitrequest & (std_2s60_burst_13_downstream_read | std_2s60_burst_13_downstream_write);
    end


  //std_2s60_burst_13_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_address != std_2s60_burst_13_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_13_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_burstcount_last_time <= std_2s60_burst_13_downstream_burstcount;
    end


  //std_2s60_burst_13_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_burstcount != std_2s60_burst_13_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_13_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_byteenable_last_time <= std_2s60_burst_13_downstream_byteenable;
    end


  //std_2s60_burst_13_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_byteenable != std_2s60_burst_13_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_13_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_read_last_time <= std_2s60_burst_13_downstream_read;
    end


  //std_2s60_burst_13_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_read != std_2s60_burst_13_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_13_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_write_last_time <= std_2s60_burst_13_downstream_write;
    end


  //std_2s60_burst_13_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_write != std_2s60_burst_13_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_13_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_13_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_13_downstream_writedata_last_time <= std_2s60_burst_13_downstream_writedata;
    end


  //std_2s60_burst_13_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_13_downstream_writedata != std_2s60_burst_13_downstream_writedata_last_time) & std_2s60_burst_13_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_13_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_14_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_14_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_14_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_14_upstream_readdata,
                                                std_2s60_burst_14_upstream_readdatavalid,
                                                std_2s60_burst_14_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_14_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_14_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_14_upstream,
                                                d1_std_2s60_burst_14_upstream_end_xfer,
                                                std_2s60_burst_14_upstream_address,
                                                std_2s60_burst_14_upstream_burstcount,
                                                std_2s60_burst_14_upstream_byteaddress,
                                                std_2s60_burst_14_upstream_byteenable,
                                                std_2s60_burst_14_upstream_debugaccess,
                                                std_2s60_burst_14_upstream_read,
                                                std_2s60_burst_14_upstream_readdata_from_sa,
                                                std_2s60_burst_14_upstream_waitrequest_from_sa,
                                                std_2s60_burst_14_upstream_write,
                                                std_2s60_burst_14_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_14_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_14_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_14_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_14_upstream;
  output           d1_std_2s60_burst_14_upstream_end_xfer;
  output  [  2: 0] std_2s60_burst_14_upstream_address;
  output  [  3: 0] std_2s60_burst_14_upstream_burstcount;
  output  [  4: 0] std_2s60_burst_14_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_14_upstream_byteenable;
  output           std_2s60_burst_14_upstream_debugaccess;
  output           std_2s60_burst_14_upstream_read;
  output  [ 31: 0] std_2s60_burst_14_upstream_readdata_from_sa;
  output           std_2s60_burst_14_upstream_waitrequest_from_sa;
  output           std_2s60_burst_14_upstream_write;
  output  [ 31: 0] std_2s60_burst_14_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_14_upstream_readdata;
  input            std_2s60_burst_14_upstream_readdatavalid;
  input            std_2s60_burst_14_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_14_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_14_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_14_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_14_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_14_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_14_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_14_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_14_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_14_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_14_upstream_from_cpu_data_master;
  wire    [  2: 0] std_2s60_burst_14_upstream_address;
  wire             std_2s60_burst_14_upstream_allgrants;
  wire             std_2s60_burst_14_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_14_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_14_upstream_any_continuerequest;
  wire             std_2s60_burst_14_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_14_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_14_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_14_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_14_upstream_bbt_burstcounter;
  wire             std_2s60_burst_14_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_14_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_14_upstream_burstcount;
  wire             std_2s60_burst_14_upstream_burstcount_fifo_empty;
  wire    [  4: 0] std_2s60_burst_14_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_14_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_14_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_14_upstream_current_burst_minus_one;
  wire             std_2s60_burst_14_upstream_debugaccess;
  wire             std_2s60_burst_14_upstream_end_xfer;
  wire             std_2s60_burst_14_upstream_firsttransfer;
  wire             std_2s60_burst_14_upstream_grant_vector;
  wire             std_2s60_burst_14_upstream_in_a_read_cycle;
  wire             std_2s60_burst_14_upstream_in_a_write_cycle;
  reg              std_2s60_burst_14_upstream_load_fifo;
  wire             std_2s60_burst_14_upstream_master_qreq_vector;
  wire             std_2s60_burst_14_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_14_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_14_upstream_next_burst_count;
  wire             std_2s60_burst_14_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_14_upstream_read;
  wire    [ 31: 0] std_2s60_burst_14_upstream_readdata_from_sa;
  wire             std_2s60_burst_14_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_14_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_14_upstream_selected_burstcount;
  reg              std_2s60_burst_14_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_14_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_14_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_14_upstream_transaction_burst_count;
  wire             std_2s60_burst_14_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_14_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_14_upstream_waits_for_read;
  wire             std_2s60_burst_14_upstream_waits_for_write;
  wire             std_2s60_burst_14_upstream_write;
  wire    [ 31: 0] std_2s60_burst_14_upstream_writedata;
  wire             wait_for_std_2s60_burst_14_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_14_upstream_end_xfer;
    end


  assign std_2s60_burst_14_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_14_upstream));
  //assign std_2s60_burst_14_upstream_readdatavalid_from_sa = std_2s60_burst_14_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_14_upstream_readdatavalid_from_sa = std_2s60_burst_14_upstream_readdatavalid;

  //assign std_2s60_burst_14_upstream_readdata_from_sa = std_2s60_burst_14_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_14_upstream_readdata_from_sa = std_2s60_burst_14_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_14_upstream = ({cpu_data_master_address_to_slave[25 : 3] , 3'b0} == 26'h2131888) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_14_upstream_waitrequest_from_sa = std_2s60_burst_14_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_14_upstream_waitrequest_from_sa = std_2s60_burst_14_upstream_waitrequest;

  //std_2s60_burst_14_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_14_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_14_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_14_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_14_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_14_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_14_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_14_upstream;

  //std_2s60_burst_14_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_14_upstream_arb_share_counter_next_value = std_2s60_burst_14_upstream_firsttransfer ? (std_2s60_burst_14_upstream_arb_share_set_values - 1) : |std_2s60_burst_14_upstream_arb_share_counter ? (std_2s60_burst_14_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_14_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_14_upstream_allgrants = |std_2s60_burst_14_upstream_grant_vector;

  //std_2s60_burst_14_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_14_upstream_end_xfer = ~(std_2s60_burst_14_upstream_waits_for_read | std_2s60_burst_14_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream = std_2s60_burst_14_upstream_end_xfer & (~std_2s60_burst_14_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_14_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_14_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream & std_2s60_burst_14_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream & ~std_2s60_burst_14_upstream_non_bursting_master_requests);

  //std_2s60_burst_14_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_14_upstream_arb_counter_enable)
          std_2s60_burst_14_upstream_arb_share_counter <= std_2s60_burst_14_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_14_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_14_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_14_upstream & ~std_2s60_burst_14_upstream_non_bursting_master_requests))
          std_2s60_burst_14_upstream_slavearbiterlockenable <= |std_2s60_burst_14_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_14/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_14_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_14_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_14_upstream_slavearbiterlockenable2 = |std_2s60_burst_14_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_14/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_14_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_14_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_14_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_14_upstream = cpu_data_master_requests_std_2s60_burst_14_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_14_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_14_upstream_move_on_to_next_transaction = std_2s60_burst_14_upstream_this_cycle_is_the_last_burst & std_2s60_burst_14_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_14_upstream, which is an e_mux
  assign std_2s60_burst_14_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_14_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_14_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_14_upstream_module burstcount_fifo_for_std_2s60_burst_14_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_14_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_14_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_14_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_14_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read & std_2s60_burst_14_upstream_load_fifo & ~(std_2s60_burst_14_upstream_this_cycle_is_the_last_burst & std_2s60_burst_14_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_14_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_14_upstream_current_burst_minus_one = std_2s60_burst_14_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_14_upstream, which is an e_mux
  assign std_2s60_burst_14_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read) & ~std_2s60_burst_14_upstream_load_fifo))? std_2s60_burst_14_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read & std_2s60_burst_14_upstream_this_cycle_is_the_last_burst & std_2s60_burst_14_upstream_burstcount_fifo_empty))? std_2s60_burst_14_upstream_selected_burstcount :
    (std_2s60_burst_14_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_14_upstream_transaction_burst_count :
    std_2s60_burst_14_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_14_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_current_burst <= 0;
      else if (std_2s60_burst_14_upstream_readdatavalid_from_sa | (~std_2s60_burst_14_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read)))
          std_2s60_burst_14_upstream_current_burst <= std_2s60_burst_14_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_14_upstream_load_fifo = (~std_2s60_burst_14_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read) & std_2s60_burst_14_upstream_load_fifo))? 1 :
    ~std_2s60_burst_14_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read) & ~std_2s60_burst_14_upstream_load_fifo | std_2s60_burst_14_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_14_upstream_load_fifo <= p0_std_2s60_burst_14_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_14_upstream, which is an e_assign
  assign std_2s60_burst_14_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_14_upstream_current_burst_minus_one) & std_2s60_burst_14_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_14_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_14_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_14_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_14_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_14_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_14_upstream),
      .full                 (),
      .read                 (std_2s60_burst_14_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_14_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_14_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_14_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_14_upstream = std_2s60_burst_14_upstream_readdatavalid_from_sa;

  //std_2s60_burst_14_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_14_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_14/upstream, which is an e_mux
  assign std_2s60_burst_14_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_14_upstream = cpu_data_master_qualified_request_std_2s60_burst_14_upstream;

  //cpu/data_master saved-grant std_2s60_burst_14/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_14_upstream = cpu_data_master_requests_std_2s60_burst_14_upstream;

  //allow new arb cycle for std_2s60_burst_14/upstream, which is an e_assign
  assign std_2s60_burst_14_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_14_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_14_upstream_master_qreq_vector = 1;

  //std_2s60_burst_14_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_14_upstream_firsttransfer = std_2s60_burst_14_upstream_begins_xfer ? std_2s60_burst_14_upstream_unreg_firsttransfer : std_2s60_burst_14_upstream_reg_firsttransfer;

  //std_2s60_burst_14_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_14_upstream_unreg_firsttransfer = ~(std_2s60_burst_14_upstream_slavearbiterlockenable & std_2s60_burst_14_upstream_any_continuerequest);

  //std_2s60_burst_14_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_14_upstream_begins_xfer)
          std_2s60_burst_14_upstream_reg_firsttransfer <= std_2s60_burst_14_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_14_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_14_upstream_next_bbt_burstcount = ((((std_2s60_burst_14_upstream_write) && (std_2s60_burst_14_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_14_upstream_burstcount - 1) :
    ((((std_2s60_burst_14_upstream_read) && (std_2s60_burst_14_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_14_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_14_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_14_upstream_begins_xfer)
          std_2s60_burst_14_upstream_bbt_burstcounter <= std_2s60_burst_14_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_14_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_14_upstream_beginbursttransfer_internal = std_2s60_burst_14_upstream_begins_xfer & (std_2s60_burst_14_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_14_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_14_upstream_read = cpu_data_master_granted_std_2s60_burst_14_upstream & cpu_data_master_read;

  //std_2s60_burst_14_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_14_upstream_write = cpu_data_master_granted_std_2s60_burst_14_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_14_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_14_upstream_address mux, which is an e_mux
  assign std_2s60_burst_14_upstream_address = shifted_address_to_std_2s60_burst_14_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_14_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_14_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_14_upstream_end_xfer <= std_2s60_burst_14_upstream_end_xfer;
    end


  //std_2s60_burst_14_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_14_upstream_waits_for_read = std_2s60_burst_14_upstream_in_a_read_cycle & std_2s60_burst_14_upstream_waitrequest_from_sa;

  //std_2s60_burst_14_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_14_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_14_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_14_upstream_in_a_read_cycle;

  //std_2s60_burst_14_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_14_upstream_waits_for_write = std_2s60_burst_14_upstream_in_a_write_cycle & std_2s60_burst_14_upstream_waitrequest_from_sa;

  //std_2s60_burst_14_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_14_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_14_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_14_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_14_upstream_counter = 0;
  //std_2s60_burst_14_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_14_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_14_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_14_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_14_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_14_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_14_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_14/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_14_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_14/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_14_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_sysid_control_slave_end_xfer,
                                                  reset_n,
                                                  std_2s60_burst_14_downstream_address,
                                                  std_2s60_burst_14_downstream_burstcount,
                                                  std_2s60_burst_14_downstream_byteenable,
                                                  std_2s60_burst_14_downstream_granted_sysid_control_slave,
                                                  std_2s60_burst_14_downstream_qualified_request_sysid_control_slave,
                                                  std_2s60_burst_14_downstream_read,
                                                  std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave,
                                                  std_2s60_burst_14_downstream_requests_sysid_control_slave,
                                                  std_2s60_burst_14_downstream_write,
                                                  std_2s60_burst_14_downstream_writedata,
                                                  sysid_control_slave_readdata_from_sa,

                                                 // outputs:
                                                  std_2s60_burst_14_downstream_address_to_slave,
                                                  std_2s60_burst_14_downstream_latency_counter,
                                                  std_2s60_burst_14_downstream_readdata,
                                                  std_2s60_burst_14_downstream_readdatavalid,
                                                  std_2s60_burst_14_downstream_reset_n,
                                                  std_2s60_burst_14_downstream_waitrequest
                                               )
;

  output  [  2: 0] std_2s60_burst_14_downstream_address_to_slave;
  output           std_2s60_burst_14_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_14_downstream_readdata;
  output           std_2s60_burst_14_downstream_readdatavalid;
  output           std_2s60_burst_14_downstream_reset_n;
  output           std_2s60_burst_14_downstream_waitrequest;
  input            clk;
  input            d1_sysid_control_slave_end_xfer;
  input            reset_n;
  input   [  2: 0] std_2s60_burst_14_downstream_address;
  input            std_2s60_burst_14_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_14_downstream_byteenable;
  input            std_2s60_burst_14_downstream_granted_sysid_control_slave;
  input            std_2s60_burst_14_downstream_qualified_request_sysid_control_slave;
  input            std_2s60_burst_14_downstream_read;
  input            std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave;
  input            std_2s60_burst_14_downstream_requests_sysid_control_slave;
  input            std_2s60_burst_14_downstream_write;
  input   [ 31: 0] std_2s60_burst_14_downstream_writedata;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  wire             pre_flush_std_2s60_burst_14_downstream_readdatavalid;
  wire             r_2;
  reg     [  2: 0] std_2s60_burst_14_downstream_address_last_time;
  wire    [  2: 0] std_2s60_burst_14_downstream_address_to_slave;
  reg              std_2s60_burst_14_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_14_downstream_byteenable_last_time;
  wire             std_2s60_burst_14_downstream_latency_counter;
  reg              std_2s60_burst_14_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_14_downstream_readdata;
  wire             std_2s60_burst_14_downstream_readdatavalid;
  wire             std_2s60_burst_14_downstream_reset_n;
  wire             std_2s60_burst_14_downstream_run;
  wire             std_2s60_burst_14_downstream_waitrequest;
  reg              std_2s60_burst_14_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_14_downstream_writedata_last_time;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (std_2s60_burst_14_downstream_qualified_request_sysid_control_slave | ~std_2s60_burst_14_downstream_requests_sysid_control_slave) & ((~std_2s60_burst_14_downstream_qualified_request_sysid_control_slave | ~std_2s60_burst_14_downstream_read | (1 & ~d1_sysid_control_slave_end_xfer & std_2s60_burst_14_downstream_read))) & ((~std_2s60_burst_14_downstream_qualified_request_sysid_control_slave | ~std_2s60_burst_14_downstream_write | (1 & std_2s60_burst_14_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_14_downstream_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_14_downstream_address_to_slave = std_2s60_burst_14_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_14_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_14_downstream_readdatavalid = 0 |
    pre_flush_std_2s60_burst_14_downstream_readdatavalid |
    std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave;

  //std_2s60_burst_14/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_14_downstream_readdata = sysid_control_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_14_downstream_waitrequest = ~std_2s60_burst_14_downstream_run;

  //latent max counter, which is an e_assign
  assign std_2s60_burst_14_downstream_latency_counter = 0;

  //std_2s60_burst_14_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_14_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_14_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_address_last_time <= std_2s60_burst_14_downstream_address;
    end


  //std_2s60_burst_14/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_14_downstream_waitrequest & (std_2s60_burst_14_downstream_read | std_2s60_burst_14_downstream_write);
    end


  //std_2s60_burst_14_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_address != std_2s60_burst_14_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_14_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_burstcount_last_time <= std_2s60_burst_14_downstream_burstcount;
    end


  //std_2s60_burst_14_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_burstcount != std_2s60_burst_14_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_14_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_byteenable_last_time <= std_2s60_burst_14_downstream_byteenable;
    end


  //std_2s60_burst_14_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_byteenable != std_2s60_burst_14_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_14_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_read_last_time <= std_2s60_burst_14_downstream_read;
    end


  //std_2s60_burst_14_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_read != std_2s60_burst_14_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_14_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_write_last_time <= std_2s60_burst_14_downstream_write;
    end


  //std_2s60_burst_14_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_write != std_2s60_burst_14_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_14_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_14_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_14_downstream_writedata_last_time <= std_2s60_burst_14_downstream_writedata;
    end


  //std_2s60_burst_14_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_14_downstream_writedata != std_2s60_burst_14_downstream_writedata_last_time) & std_2s60_burst_14_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_14_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_15_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  wire             full_9;
  reg     [  4: 0] how_many_ones;
  wire    [  4: 0] one_count_minus_one;
  wire    [  4: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_8;
  wire    [  4: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_8;
  assign empty = !full_0;
  assign full_9 = 0;
  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    0;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_15_upstream_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  wire             full_9;
  reg     [  4: 0] how_many_ones;
  wire    [  4: 0] one_count_minus_one;
  wire    [  4: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  wire    [  4: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_8;
  assign empty = !full_0;
  assign full_9 = 0;
  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    0;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_15_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_instruction_master_address_to_slave,
                                                cpu_instruction_master_burstcount,
                                                cpu_instruction_master_latency_counter,
                                                cpu_instruction_master_read,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                                reset_n,
                                                std_2s60_burst_15_upstream_readdata,
                                                std_2s60_burst_15_upstream_readdatavalid,
                                                std_2s60_burst_15_upstream_waitrequest,

                                               // outputs:
                                                cpu_instruction_master_granted_std_2s60_burst_15_upstream,
                                                cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                                cpu_instruction_master_requests_std_2s60_burst_15_upstream,
                                                d1_std_2s60_burst_15_upstream_end_xfer,
                                                std_2s60_burst_15_upstream_address,
                                                std_2s60_burst_15_upstream_byteaddress,
                                                std_2s60_burst_15_upstream_byteenable,
                                                std_2s60_burst_15_upstream_debugaccess,
                                                std_2s60_burst_15_upstream_read,
                                                std_2s60_burst_15_upstream_readdata_from_sa,
                                                std_2s60_burst_15_upstream_waitrequest_from_sa,
                                                std_2s60_burst_15_upstream_write
                                             )
;

  output           cpu_instruction_master_granted_std_2s60_burst_15_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_15_upstream;
  output           d1_std_2s60_burst_15_upstream_end_xfer;
  output  [ 23: 0] std_2s60_burst_15_upstream_address;
  output  [ 25: 0] std_2s60_burst_15_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_15_upstream_byteenable;
  output           std_2s60_burst_15_upstream_debugaccess;
  output           std_2s60_burst_15_upstream_read;
  output  [ 31: 0] std_2s60_burst_15_upstream_readdata_from_sa;
  output           std_2s60_burst_15_upstream_waitrequest_from_sa;
  output           std_2s60_burst_15_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_15_upstream_readdata;
  input            std_2s60_burst_15_upstream_readdatavalid;
  input            std_2s60_burst_15_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_15_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_15_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_15_upstream_load_fifo;
  wire    [ 23: 0] std_2s60_burst_15_upstream_address;
  wire             std_2s60_burst_15_upstream_allgrants;
  wire             std_2s60_burst_15_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_15_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_15_upstream_any_continuerequest;
  wire             std_2s60_burst_15_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_15_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_15_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_15_upstream_arb_share_set_values;
  wire             std_2s60_burst_15_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_15_upstream_begins_xfer;
  wire             std_2s60_burst_15_upstream_burstcount_fifo_empty;
  wire    [ 25: 0] std_2s60_burst_15_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_15_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_15_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_15_upstream_current_burst_minus_one;
  wire             std_2s60_burst_15_upstream_debugaccess;
  wire             std_2s60_burst_15_upstream_end_xfer;
  wire             std_2s60_burst_15_upstream_firsttransfer;
  wire             std_2s60_burst_15_upstream_grant_vector;
  wire             std_2s60_burst_15_upstream_in_a_read_cycle;
  wire             std_2s60_burst_15_upstream_in_a_write_cycle;
  reg              std_2s60_burst_15_upstream_load_fifo;
  wire             std_2s60_burst_15_upstream_master_qreq_vector;
  wire             std_2s60_burst_15_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_15_upstream_next_burst_count;
  wire             std_2s60_burst_15_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_15_upstream_read;
  wire    [ 31: 0] std_2s60_burst_15_upstream_readdata_from_sa;
  wire             std_2s60_burst_15_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_15_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_15_upstream_selected_burstcount;
  reg              std_2s60_burst_15_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_15_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_15_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_15_upstream_transaction_burst_count;
  wire             std_2s60_burst_15_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_15_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_15_upstream_waits_for_read;
  wire             std_2s60_burst_15_upstream_waits_for_write;
  wire             std_2s60_burst_15_upstream_write;
  wire             wait_for_std_2s60_burst_15_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_15_upstream_end_xfer;
    end


  assign std_2s60_burst_15_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream));
  //assign std_2s60_burst_15_upstream_readdatavalid_from_sa = std_2s60_burst_15_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_15_upstream_readdatavalid_from_sa = std_2s60_burst_15_upstream_readdatavalid;

  //assign std_2s60_burst_15_upstream_readdata_from_sa = std_2s60_burst_15_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_15_upstream_readdata_from_sa = std_2s60_burst_15_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_15_upstream = (({cpu_instruction_master_address_to_slave[25 : 24] , 24'b0} == 26'h1000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_15_upstream_waitrequest_from_sa = std_2s60_burst_15_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_15_upstream_waitrequest_from_sa = std_2s60_burst_15_upstream_waitrequest;

  //std_2s60_burst_15_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_15_upstream_arb_share_set_values = 1;

  //std_2s60_burst_15_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_15_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_15_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_15_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_15_upstream;

  //std_2s60_burst_15_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_15_upstream_arb_share_counter_next_value = std_2s60_burst_15_upstream_firsttransfer ? (std_2s60_burst_15_upstream_arb_share_set_values - 1) : |std_2s60_burst_15_upstream_arb_share_counter ? (std_2s60_burst_15_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_15_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_15_upstream_allgrants = |std_2s60_burst_15_upstream_grant_vector;

  //std_2s60_burst_15_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_15_upstream_end_xfer = ~(std_2s60_burst_15_upstream_waits_for_read | std_2s60_burst_15_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream = std_2s60_burst_15_upstream_end_xfer & (~std_2s60_burst_15_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_15_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_15_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream & std_2s60_burst_15_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream & ~std_2s60_burst_15_upstream_non_bursting_master_requests);

  //std_2s60_burst_15_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_15_upstream_arb_counter_enable)
          std_2s60_burst_15_upstream_arb_share_counter <= std_2s60_burst_15_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_15_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_15_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_15_upstream & ~std_2s60_burst_15_upstream_non_bursting_master_requests))
          std_2s60_burst_15_upstream_slavearbiterlockenable <= |std_2s60_burst_15_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_15/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_15_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_15_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_15_upstream_slavearbiterlockenable2 = |std_2s60_burst_15_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_15/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_15_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_15_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_15_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream = cpu_instruction_master_requests_std_2s60_burst_15_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_15_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_15_upstream_move_on_to_next_transaction = std_2s60_burst_15_upstream_this_cycle_is_the_last_burst & std_2s60_burst_15_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_15_upstream, which is an e_mux
  assign std_2s60_burst_15_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_15_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_15_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_15_upstream_module burstcount_fifo_for_std_2s60_burst_15_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_15_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_15_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_15_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_15_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read & std_2s60_burst_15_upstream_load_fifo & ~(std_2s60_burst_15_upstream_this_cycle_is_the_last_burst & std_2s60_burst_15_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_15_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_15_upstream_current_burst_minus_one = std_2s60_burst_15_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_15_upstream, which is an e_mux
  assign std_2s60_burst_15_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read) & ~std_2s60_burst_15_upstream_load_fifo))? std_2s60_burst_15_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read & std_2s60_burst_15_upstream_this_cycle_is_the_last_burst & std_2s60_burst_15_upstream_burstcount_fifo_empty))? std_2s60_burst_15_upstream_selected_burstcount :
    (std_2s60_burst_15_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_15_upstream_transaction_burst_count :
    std_2s60_burst_15_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_15_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_upstream_current_burst <= 0;
      else if (std_2s60_burst_15_upstream_readdatavalid_from_sa | (~std_2s60_burst_15_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read)))
          std_2s60_burst_15_upstream_current_burst <= std_2s60_burst_15_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_15_upstream_load_fifo = (~std_2s60_burst_15_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read) & std_2s60_burst_15_upstream_load_fifo))? 1 :
    ~std_2s60_burst_15_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read) & ~std_2s60_burst_15_upstream_load_fifo | std_2s60_burst_15_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_15_upstream_load_fifo <= p0_std_2s60_burst_15_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_15_upstream, which is an e_assign
  assign std_2s60_burst_15_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_15_upstream_current_burst_minus_one) & std_2s60_burst_15_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_15_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_15_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_15_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_15_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_15_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_15_upstream),
      .full                 (),
      .read                 (std_2s60_burst_15_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_15_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_15_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream = std_2s60_burst_15_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_15/upstream, which is an e_mux
  assign std_2s60_burst_15_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_15_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_15/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_15_upstream = cpu_instruction_master_requests_std_2s60_burst_15_upstream;

  //allow new arb cycle for std_2s60_burst_15/upstream, which is an e_assign
  assign std_2s60_burst_15_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_15_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_15_upstream_master_qreq_vector = 1;

  //std_2s60_burst_15_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_15_upstream_firsttransfer = std_2s60_burst_15_upstream_begins_xfer ? std_2s60_burst_15_upstream_unreg_firsttransfer : std_2s60_burst_15_upstream_reg_firsttransfer;

  //std_2s60_burst_15_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_15_upstream_unreg_firsttransfer = ~(std_2s60_burst_15_upstream_slavearbiterlockenable & std_2s60_burst_15_upstream_any_continuerequest);

  //std_2s60_burst_15_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_15_upstream_begins_xfer)
          std_2s60_burst_15_upstream_reg_firsttransfer <= std_2s60_burst_15_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_15_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_15_upstream_beginbursttransfer_internal = std_2s60_burst_15_upstream_begins_xfer;

  //std_2s60_burst_15_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_15_upstream_read = cpu_instruction_master_granted_std_2s60_burst_15_upstream & cpu_instruction_master_read;

  //std_2s60_burst_15_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_15_upstream_write = 0;

  //std_2s60_burst_15_upstream_address mux, which is an e_mux
  assign std_2s60_burst_15_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_std_2s60_burst_15_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_15_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_15_upstream_end_xfer <= std_2s60_burst_15_upstream_end_xfer;
    end


  //std_2s60_burst_15_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_15_upstream_waits_for_read = std_2s60_burst_15_upstream_in_a_read_cycle & std_2s60_burst_15_upstream_waitrequest_from_sa;

  //std_2s60_burst_15_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_15_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_15_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_15_upstream_in_a_read_cycle;

  //std_2s60_burst_15_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_15_upstream_waits_for_write = std_2s60_burst_15_upstream_in_a_write_cycle & std_2s60_burst_15_upstream_waitrequest_from_sa;

  //std_2s60_burst_15_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_15_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_15_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_15_upstream_counter = 0;
  //std_2s60_burst_15_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_15_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_15_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_15/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_15_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_15/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_15_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_sdram_s1_end_xfer,
                                                  reset_n,
                                                  sdram_s1_readdata_from_sa,
                                                  sdram_s1_waitrequest_from_sa,
                                                  std_2s60_burst_15_downstream_address,
                                                  std_2s60_burst_15_downstream_burstcount,
                                                  std_2s60_burst_15_downstream_byteenable,
                                                  std_2s60_burst_15_downstream_granted_sdram_s1,
                                                  std_2s60_burst_15_downstream_qualified_request_sdram_s1,
                                                  std_2s60_burst_15_downstream_read,
                                                  std_2s60_burst_15_downstream_read_data_valid_sdram_s1,
                                                  std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register,
                                                  std_2s60_burst_15_downstream_requests_sdram_s1,
                                                  std_2s60_burst_15_downstream_write,
                                                  std_2s60_burst_15_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_15_downstream_address_to_slave,
                                                  std_2s60_burst_15_downstream_latency_counter,
                                                  std_2s60_burst_15_downstream_readdata,
                                                  std_2s60_burst_15_downstream_readdatavalid,
                                                  std_2s60_burst_15_downstream_reset_n,
                                                  std_2s60_burst_15_downstream_waitrequest
                                               )
;

  output  [ 23: 0] std_2s60_burst_15_downstream_address_to_slave;
  output           std_2s60_burst_15_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_15_downstream_readdata;
  output           std_2s60_burst_15_downstream_readdatavalid;
  output           std_2s60_burst_15_downstream_reset_n;
  output           std_2s60_burst_15_downstream_waitrequest;
  input            clk;
  input            d1_sdram_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sdram_s1_readdata_from_sa;
  input            sdram_s1_waitrequest_from_sa;
  input   [ 23: 0] std_2s60_burst_15_downstream_address;
  input            std_2s60_burst_15_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_15_downstream_byteenable;
  input            std_2s60_burst_15_downstream_granted_sdram_s1;
  input            std_2s60_burst_15_downstream_qualified_request_sdram_s1;
  input            std_2s60_burst_15_downstream_read;
  input            std_2s60_burst_15_downstream_read_data_valid_sdram_s1;
  input            std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register;
  input            std_2s60_burst_15_downstream_requests_sdram_s1;
  input            std_2s60_burst_15_downstream_write;
  input   [ 31: 0] std_2s60_burst_15_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_15_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_15_downstream_readdatavalid;
  wire             r_0;
  reg     [ 23: 0] std_2s60_burst_15_downstream_address_last_time;
  wire    [ 23: 0] std_2s60_burst_15_downstream_address_to_slave;
  reg              std_2s60_burst_15_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_15_downstream_byteenable_last_time;
  wire             std_2s60_burst_15_downstream_is_granted_some_slave;
  reg              std_2s60_burst_15_downstream_latency_counter;
  reg              std_2s60_burst_15_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_15_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_15_downstream_readdata;
  wire             std_2s60_burst_15_downstream_readdatavalid;
  wire             std_2s60_burst_15_downstream_reset_n;
  wire             std_2s60_burst_15_downstream_run;
  wire             std_2s60_burst_15_downstream_waitrequest;
  reg              std_2s60_burst_15_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_15_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_15_downstream_qualified_request_sdram_s1 | ~std_2s60_burst_15_downstream_requests_sdram_s1) & (std_2s60_burst_15_downstream_granted_sdram_s1 | ~std_2s60_burst_15_downstream_qualified_request_sdram_s1) & ((~std_2s60_burst_15_downstream_qualified_request_sdram_s1 | ~(std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write) | (1 & ~sdram_s1_waitrequest_from_sa & (std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write)))) & ((~std_2s60_burst_15_downstream_qualified_request_sdram_s1 | ~(std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write) | (1 & ~sdram_s1_waitrequest_from_sa & (std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_15_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_15_downstream_address_to_slave = std_2s60_burst_15_downstream_address;

  //std_2s60_burst_15_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_15_downstream_read_but_no_slave_selected <= std_2s60_burst_15_downstream_read & std_2s60_burst_15_downstream_run & ~std_2s60_burst_15_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_15_downstream_is_granted_some_slave = std_2s60_burst_15_downstream_granted_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_15_downstream_readdatavalid = std_2s60_burst_15_downstream_read_data_valid_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_15_downstream_readdatavalid = std_2s60_burst_15_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_15_downstream_readdatavalid;

  //std_2s60_burst_15/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_15_downstream_readdata = sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_15_downstream_waitrequest = ~std_2s60_burst_15_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_15_downstream_latency_counter <= p1_std_2s60_burst_15_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_15_downstream_latency_counter = ((std_2s60_burst_15_downstream_run & std_2s60_burst_15_downstream_read))? latency_load_value :
    (std_2s60_burst_15_downstream_latency_counter)? std_2s60_burst_15_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //std_2s60_burst_15_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_15_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_15_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_address_last_time <= std_2s60_burst_15_downstream_address;
    end


  //std_2s60_burst_15/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_15_downstream_waitrequest & (std_2s60_burst_15_downstream_read | std_2s60_burst_15_downstream_write);
    end


  //std_2s60_burst_15_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_address != std_2s60_burst_15_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_15_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_burstcount_last_time <= std_2s60_burst_15_downstream_burstcount;
    end


  //std_2s60_burst_15_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_burstcount != std_2s60_burst_15_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_15_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_byteenable_last_time <= std_2s60_burst_15_downstream_byteenable;
    end


  //std_2s60_burst_15_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_byteenable != std_2s60_burst_15_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_15_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_read_last_time <= std_2s60_burst_15_downstream_read;
    end


  //std_2s60_burst_15_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_read != std_2s60_burst_15_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_15_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_write_last_time <= std_2s60_burst_15_downstream_write;
    end


  //std_2s60_burst_15_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_write != std_2s60_burst_15_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_15_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_15_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_15_downstream_writedata_last_time <= std_2s60_burst_15_downstream_writedata;
    end


  //std_2s60_burst_15_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_15_downstream_writedata != std_2s60_burst_15_downstream_writedata_last_time) & std_2s60_burst_15_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_15_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_16_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  wire             full_9;
  reg     [  4: 0] how_many_ones;
  wire    [  4: 0] one_count_minus_one;
  wire    [  4: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_8;
  wire    [  4: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_8;
  assign empty = !full_0;
  assign full_9 = 0;
  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    0;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_16_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  wire             full_9;
  reg     [  4: 0] how_many_ones;
  wire    [  4: 0] one_count_minus_one;
  wire    [  4: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  wire    [  4: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_8;
  assign empty = !full_0;
  assign full_9 = 0;
  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    0;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_16_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_16_upstream_readdata,
                                                std_2s60_burst_16_upstream_readdatavalid,
                                                std_2s60_burst_16_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_16_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_16_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_16_upstream,
                                                d1_std_2s60_burst_16_upstream_end_xfer,
                                                std_2s60_burst_16_upstream_address,
                                                std_2s60_burst_16_upstream_burstcount,
                                                std_2s60_burst_16_upstream_byteaddress,
                                                std_2s60_burst_16_upstream_byteenable,
                                                std_2s60_burst_16_upstream_debugaccess,
                                                std_2s60_burst_16_upstream_read,
                                                std_2s60_burst_16_upstream_readdata_from_sa,
                                                std_2s60_burst_16_upstream_waitrequest_from_sa,
                                                std_2s60_burst_16_upstream_write,
                                                std_2s60_burst_16_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_16_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_16_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_16_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_16_upstream;
  output           d1_std_2s60_burst_16_upstream_end_xfer;
  output  [ 23: 0] std_2s60_burst_16_upstream_address;
  output  [  3: 0] std_2s60_burst_16_upstream_burstcount;
  output  [ 25: 0] std_2s60_burst_16_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_16_upstream_byteenable;
  output           std_2s60_burst_16_upstream_debugaccess;
  output           std_2s60_burst_16_upstream_read;
  output  [ 31: 0] std_2s60_burst_16_upstream_readdata_from_sa;
  output           std_2s60_burst_16_upstream_waitrequest_from_sa;
  output           std_2s60_burst_16_upstream_write;
  output  [ 31: 0] std_2s60_burst_16_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_16_upstream_readdata;
  input            std_2s60_burst_16_upstream_readdatavalid;
  input            std_2s60_burst_16_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_16_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_16_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_16_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_16_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_16_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_16_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_16_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_16_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_16_upstream_load_fifo;
  wire    [ 23: 0] std_2s60_burst_16_upstream_address;
  wire             std_2s60_burst_16_upstream_allgrants;
  wire             std_2s60_burst_16_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_16_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_16_upstream_any_continuerequest;
  wire             std_2s60_burst_16_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_16_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_16_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_16_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_16_upstream_bbt_burstcounter;
  wire             std_2s60_burst_16_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_16_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_16_upstream_burstcount;
  wire             std_2s60_burst_16_upstream_burstcount_fifo_empty;
  wire    [ 25: 0] std_2s60_burst_16_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_16_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_16_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_16_upstream_current_burst_minus_one;
  wire             std_2s60_burst_16_upstream_debugaccess;
  wire             std_2s60_burst_16_upstream_end_xfer;
  wire             std_2s60_burst_16_upstream_firsttransfer;
  wire             std_2s60_burst_16_upstream_grant_vector;
  wire             std_2s60_burst_16_upstream_in_a_read_cycle;
  wire             std_2s60_burst_16_upstream_in_a_write_cycle;
  reg              std_2s60_burst_16_upstream_load_fifo;
  wire             std_2s60_burst_16_upstream_master_qreq_vector;
  wire             std_2s60_burst_16_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_16_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_16_upstream_next_burst_count;
  wire             std_2s60_burst_16_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_16_upstream_read;
  wire    [ 31: 0] std_2s60_burst_16_upstream_readdata_from_sa;
  wire             std_2s60_burst_16_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_16_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_16_upstream_selected_burstcount;
  reg              std_2s60_burst_16_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_16_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_16_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_16_upstream_transaction_burst_count;
  wire             std_2s60_burst_16_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_16_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_16_upstream_waits_for_read;
  wire             std_2s60_burst_16_upstream_waits_for_write;
  wire             std_2s60_burst_16_upstream_write;
  wire    [ 31: 0] std_2s60_burst_16_upstream_writedata;
  wire             wait_for_std_2s60_burst_16_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_16_upstream_end_xfer;
    end


  assign std_2s60_burst_16_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_16_upstream));
  //assign std_2s60_burst_16_upstream_readdatavalid_from_sa = std_2s60_burst_16_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_16_upstream_readdatavalid_from_sa = std_2s60_burst_16_upstream_readdatavalid;

  //assign std_2s60_burst_16_upstream_readdata_from_sa = std_2s60_burst_16_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_16_upstream_readdata_from_sa = std_2s60_burst_16_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_16_upstream = ({cpu_data_master_address_to_slave[25 : 24] , 24'b0} == 26'h1000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_16_upstream_waitrequest_from_sa = std_2s60_burst_16_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_16_upstream_waitrequest_from_sa = std_2s60_burst_16_upstream_waitrequest;

  //std_2s60_burst_16_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_16_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_16_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_16_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_16_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_16_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_16_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_16_upstream;

  //std_2s60_burst_16_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_16_upstream_arb_share_counter_next_value = std_2s60_burst_16_upstream_firsttransfer ? (std_2s60_burst_16_upstream_arb_share_set_values - 1) : |std_2s60_burst_16_upstream_arb_share_counter ? (std_2s60_burst_16_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_16_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_16_upstream_allgrants = |std_2s60_burst_16_upstream_grant_vector;

  //std_2s60_burst_16_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_16_upstream_end_xfer = ~(std_2s60_burst_16_upstream_waits_for_read | std_2s60_burst_16_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream = std_2s60_burst_16_upstream_end_xfer & (~std_2s60_burst_16_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_16_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_16_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream & std_2s60_burst_16_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream & ~std_2s60_burst_16_upstream_non_bursting_master_requests);

  //std_2s60_burst_16_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_16_upstream_arb_counter_enable)
          std_2s60_burst_16_upstream_arb_share_counter <= std_2s60_burst_16_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_16_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_16_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_16_upstream & ~std_2s60_burst_16_upstream_non_bursting_master_requests))
          std_2s60_burst_16_upstream_slavearbiterlockenable <= |std_2s60_burst_16_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_16/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_16_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_16_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_16_upstream_slavearbiterlockenable2 = |std_2s60_burst_16_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_16/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_16_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_16_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_16_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_16_upstream = cpu_data_master_requests_std_2s60_burst_16_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_16_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_16_upstream_move_on_to_next_transaction = std_2s60_burst_16_upstream_this_cycle_is_the_last_burst & std_2s60_burst_16_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_16_upstream, which is an e_mux
  assign std_2s60_burst_16_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_16_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_16_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_16_upstream_module burstcount_fifo_for_std_2s60_burst_16_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_16_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_16_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_16_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_16_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read & std_2s60_burst_16_upstream_load_fifo & ~(std_2s60_burst_16_upstream_this_cycle_is_the_last_burst & std_2s60_burst_16_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_16_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_16_upstream_current_burst_minus_one = std_2s60_burst_16_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_16_upstream, which is an e_mux
  assign std_2s60_burst_16_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read) & ~std_2s60_burst_16_upstream_load_fifo))? std_2s60_burst_16_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read & std_2s60_burst_16_upstream_this_cycle_is_the_last_burst & std_2s60_burst_16_upstream_burstcount_fifo_empty))? std_2s60_burst_16_upstream_selected_burstcount :
    (std_2s60_burst_16_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_16_upstream_transaction_burst_count :
    std_2s60_burst_16_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_16_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_current_burst <= 0;
      else if (std_2s60_burst_16_upstream_readdatavalid_from_sa | (~std_2s60_burst_16_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read)))
          std_2s60_burst_16_upstream_current_burst <= std_2s60_burst_16_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_16_upstream_load_fifo = (~std_2s60_burst_16_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read) & std_2s60_burst_16_upstream_load_fifo))? 1 :
    ~std_2s60_burst_16_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read) & ~std_2s60_burst_16_upstream_load_fifo | std_2s60_burst_16_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_16_upstream_load_fifo <= p0_std_2s60_burst_16_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_16_upstream, which is an e_assign
  assign std_2s60_burst_16_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_16_upstream_current_burst_minus_one) & std_2s60_burst_16_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_16_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_16_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_16_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_16_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_16_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_16_upstream),
      .full                 (),
      .read                 (std_2s60_burst_16_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_16_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_16_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_16_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_16_upstream = std_2s60_burst_16_upstream_readdatavalid_from_sa;

  //std_2s60_burst_16_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_16_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_16/upstream, which is an e_mux
  assign std_2s60_burst_16_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_16_upstream = cpu_data_master_qualified_request_std_2s60_burst_16_upstream;

  //cpu/data_master saved-grant std_2s60_burst_16/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_16_upstream = cpu_data_master_requests_std_2s60_burst_16_upstream;

  //allow new arb cycle for std_2s60_burst_16/upstream, which is an e_assign
  assign std_2s60_burst_16_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_16_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_16_upstream_master_qreq_vector = 1;

  //std_2s60_burst_16_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_16_upstream_firsttransfer = std_2s60_burst_16_upstream_begins_xfer ? std_2s60_burst_16_upstream_unreg_firsttransfer : std_2s60_burst_16_upstream_reg_firsttransfer;

  //std_2s60_burst_16_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_16_upstream_unreg_firsttransfer = ~(std_2s60_burst_16_upstream_slavearbiterlockenable & std_2s60_burst_16_upstream_any_continuerequest);

  //std_2s60_burst_16_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_16_upstream_begins_xfer)
          std_2s60_burst_16_upstream_reg_firsttransfer <= std_2s60_burst_16_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_16_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_16_upstream_next_bbt_burstcount = ((((std_2s60_burst_16_upstream_write) && (std_2s60_burst_16_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_16_upstream_burstcount - 1) :
    ((((std_2s60_burst_16_upstream_read) && (std_2s60_burst_16_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_16_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_16_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_16_upstream_begins_xfer)
          std_2s60_burst_16_upstream_bbt_burstcounter <= std_2s60_burst_16_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_16_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_16_upstream_beginbursttransfer_internal = std_2s60_burst_16_upstream_begins_xfer & (std_2s60_burst_16_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_16_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_16_upstream_read = cpu_data_master_granted_std_2s60_burst_16_upstream & cpu_data_master_read;

  //std_2s60_burst_16_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_16_upstream_write = cpu_data_master_granted_std_2s60_burst_16_upstream & cpu_data_master_write;

  //std_2s60_burst_16_upstream_address mux, which is an e_mux
  assign std_2s60_burst_16_upstream_address = cpu_data_master_address_to_slave;

  //d1_std_2s60_burst_16_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_16_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_16_upstream_end_xfer <= std_2s60_burst_16_upstream_end_xfer;
    end


  //std_2s60_burst_16_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_16_upstream_waits_for_read = std_2s60_burst_16_upstream_in_a_read_cycle & std_2s60_burst_16_upstream_waitrequest_from_sa;

  //std_2s60_burst_16_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_16_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_16_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_16_upstream_in_a_read_cycle;

  //std_2s60_burst_16_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_16_upstream_waits_for_write = std_2s60_burst_16_upstream_in_a_write_cycle & std_2s60_burst_16_upstream_waitrequest_from_sa;

  //std_2s60_burst_16_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_16_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_16_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_16_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_16_upstream_counter = 0;
  //std_2s60_burst_16_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_16_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_16_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_16_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_16_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_16_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_16_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_16/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_16_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_16/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_16_downstream_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  d1_sdram_s1_end_xfer,
                                                  reset_n,
                                                  sdram_s1_readdata_from_sa,
                                                  sdram_s1_waitrequest_from_sa,
                                                  std_2s60_burst_16_downstream_address,
                                                  std_2s60_burst_16_downstream_burstcount,
                                                  std_2s60_burst_16_downstream_byteenable,
                                                  std_2s60_burst_16_downstream_granted_sdram_s1,
                                                  std_2s60_burst_16_downstream_qualified_request_sdram_s1,
                                                  std_2s60_burst_16_downstream_read,
                                                  std_2s60_burst_16_downstream_read_data_valid_sdram_s1,
                                                  std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register,
                                                  std_2s60_burst_16_downstream_requests_sdram_s1,
                                                  std_2s60_burst_16_downstream_write,
                                                  std_2s60_burst_16_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_16_downstream_address_to_slave,
                                                  std_2s60_burst_16_downstream_latency_counter,
                                                  std_2s60_burst_16_downstream_readdata,
                                                  std_2s60_burst_16_downstream_readdatavalid,
                                                  std_2s60_burst_16_downstream_reset_n,
                                                  std_2s60_burst_16_downstream_waitrequest
                                               )
;

  output  [ 23: 0] std_2s60_burst_16_downstream_address_to_slave;
  output           std_2s60_burst_16_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_16_downstream_readdata;
  output           std_2s60_burst_16_downstream_readdatavalid;
  output           std_2s60_burst_16_downstream_reset_n;
  output           std_2s60_burst_16_downstream_waitrequest;
  input            clk;
  input            d1_sdram_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sdram_s1_readdata_from_sa;
  input            sdram_s1_waitrequest_from_sa;
  input   [ 23: 0] std_2s60_burst_16_downstream_address;
  input            std_2s60_burst_16_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_16_downstream_byteenable;
  input            std_2s60_burst_16_downstream_granted_sdram_s1;
  input            std_2s60_burst_16_downstream_qualified_request_sdram_s1;
  input            std_2s60_burst_16_downstream_read;
  input            std_2s60_burst_16_downstream_read_data_valid_sdram_s1;
  input            std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register;
  input            std_2s60_burst_16_downstream_requests_sdram_s1;
  input            std_2s60_burst_16_downstream_write;
  input   [ 31: 0] std_2s60_burst_16_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_16_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_16_downstream_readdatavalid;
  wire             r_0;
  reg     [ 23: 0] std_2s60_burst_16_downstream_address_last_time;
  wire    [ 23: 0] std_2s60_burst_16_downstream_address_to_slave;
  reg              std_2s60_burst_16_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_16_downstream_byteenable_last_time;
  wire             std_2s60_burst_16_downstream_is_granted_some_slave;
  reg              std_2s60_burst_16_downstream_latency_counter;
  reg              std_2s60_burst_16_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_16_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_16_downstream_readdata;
  wire             std_2s60_burst_16_downstream_readdatavalid;
  wire             std_2s60_burst_16_downstream_reset_n;
  wire             std_2s60_burst_16_downstream_run;
  wire             std_2s60_burst_16_downstream_waitrequest;
  reg              std_2s60_burst_16_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_16_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_16_downstream_qualified_request_sdram_s1 | ~std_2s60_burst_16_downstream_requests_sdram_s1) & (std_2s60_burst_16_downstream_granted_sdram_s1 | ~std_2s60_burst_16_downstream_qualified_request_sdram_s1) & ((~std_2s60_burst_16_downstream_qualified_request_sdram_s1 | ~(std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write) | (1 & ~sdram_s1_waitrequest_from_sa & (std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write)))) & ((~std_2s60_burst_16_downstream_qualified_request_sdram_s1 | ~(std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write) | (1 & ~sdram_s1_waitrequest_from_sa & (std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_16_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_16_downstream_address_to_slave = std_2s60_burst_16_downstream_address;

  //std_2s60_burst_16_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_16_downstream_read_but_no_slave_selected <= std_2s60_burst_16_downstream_read & std_2s60_burst_16_downstream_run & ~std_2s60_burst_16_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_16_downstream_is_granted_some_slave = std_2s60_burst_16_downstream_granted_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_16_downstream_readdatavalid = std_2s60_burst_16_downstream_read_data_valid_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_16_downstream_readdatavalid = std_2s60_burst_16_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_16_downstream_readdatavalid;

  //std_2s60_burst_16/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_16_downstream_readdata = sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_16_downstream_waitrequest = ~std_2s60_burst_16_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_16_downstream_latency_counter <= p1_std_2s60_burst_16_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_16_downstream_latency_counter = ((std_2s60_burst_16_downstream_run & std_2s60_burst_16_downstream_read))? latency_load_value :
    (std_2s60_burst_16_downstream_latency_counter)? std_2s60_burst_16_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //std_2s60_burst_16_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_16_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_16_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_address_last_time <= std_2s60_burst_16_downstream_address;
    end


  //std_2s60_burst_16/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_16_downstream_waitrequest & (std_2s60_burst_16_downstream_read | std_2s60_burst_16_downstream_write);
    end


  //std_2s60_burst_16_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_address != std_2s60_burst_16_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_16_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_burstcount_last_time <= std_2s60_burst_16_downstream_burstcount;
    end


  //std_2s60_burst_16_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_burstcount != std_2s60_burst_16_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_16_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_byteenable_last_time <= std_2s60_burst_16_downstream_byteenable;
    end


  //std_2s60_burst_16_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_byteenable != std_2s60_burst_16_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_16_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_read_last_time <= std_2s60_burst_16_downstream_read;
    end


  //std_2s60_burst_16_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_read != std_2s60_burst_16_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_16_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_write_last_time <= std_2s60_burst_16_downstream_write;
    end


  //std_2s60_burst_16_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_write != std_2s60_burst_16_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_16_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_16_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_16_downstream_writedata_last_time <= std_2s60_burst_16_downstream_writedata;
    end


  //std_2s60_burst_16_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_16_downstream_writedata != std_2s60_burst_16_downstream_writedata_last_time) & std_2s60_burst_16_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_16_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_17_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_17_upstream_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_17_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_burstcount,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_debugaccess,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                                cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,
                                                std_2s60_burst_17_upstream_readdata,
                                                std_2s60_burst_17_upstream_readdatavalid,
                                                std_2s60_burst_17_upstream_waitrequest,

                                               // outputs:
                                                cpu_data_master_granted_std_2s60_burst_17_upstream,
                                                cpu_data_master_qualified_request_std_2s60_burst_17_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream,
                                                cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                                cpu_data_master_requests_std_2s60_burst_17_upstream,
                                                d1_std_2s60_burst_17_upstream_end_xfer,
                                                std_2s60_burst_17_upstream_address,
                                                std_2s60_burst_17_upstream_burstcount,
                                                std_2s60_burst_17_upstream_byteaddress,
                                                std_2s60_burst_17_upstream_byteenable,
                                                std_2s60_burst_17_upstream_debugaccess,
                                                std_2s60_burst_17_upstream_read,
                                                std_2s60_burst_17_upstream_readdata_from_sa,
                                                std_2s60_burst_17_upstream_waitrequest_from_sa,
                                                std_2s60_burst_17_upstream_write,
                                                std_2s60_burst_17_upstream_writedata
                                             )
;

  output           cpu_data_master_granted_std_2s60_burst_17_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_17_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_17_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_17_upstream;
  output           d1_std_2s60_burst_17_upstream_end_xfer;
  output  [ 13: 0] std_2s60_burst_17_upstream_address;
  output  [  3: 0] std_2s60_burst_17_upstream_burstcount;
  output  [ 15: 0] std_2s60_burst_17_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_17_upstream_byteenable;
  output           std_2s60_burst_17_upstream_debugaccess;
  output           std_2s60_burst_17_upstream_read;
  output  [ 31: 0] std_2s60_burst_17_upstream_readdata_from_sa;
  output           std_2s60_burst_17_upstream_waitrequest_from_sa;
  output           std_2s60_burst_17_upstream_write;
  output  [ 31: 0] std_2s60_burst_17_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_17_upstream_readdata;
  input            std_2s60_burst_17_upstream_readdatavalid;
  input            std_2s60_burst_17_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_17_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_17_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_17_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_17_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_17_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_17_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_17_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_17_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_17_upstream_load_fifo;
  wire    [ 13: 0] std_2s60_burst_17_upstream_address;
  wire             std_2s60_burst_17_upstream_allgrants;
  wire             std_2s60_burst_17_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_17_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_17_upstream_any_continuerequest;
  wire             std_2s60_burst_17_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_17_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_17_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_17_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_17_upstream_bbt_burstcounter;
  wire             std_2s60_burst_17_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_17_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_17_upstream_burstcount;
  wire             std_2s60_burst_17_upstream_burstcount_fifo_empty;
  wire    [ 15: 0] std_2s60_burst_17_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_17_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_17_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_17_upstream_current_burst_minus_one;
  wire             std_2s60_burst_17_upstream_debugaccess;
  wire             std_2s60_burst_17_upstream_end_xfer;
  wire             std_2s60_burst_17_upstream_firsttransfer;
  wire             std_2s60_burst_17_upstream_grant_vector;
  wire             std_2s60_burst_17_upstream_in_a_read_cycle;
  wire             std_2s60_burst_17_upstream_in_a_write_cycle;
  reg              std_2s60_burst_17_upstream_load_fifo;
  wire             std_2s60_burst_17_upstream_master_qreq_vector;
  wire             std_2s60_burst_17_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_17_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_17_upstream_next_burst_count;
  wire             std_2s60_burst_17_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_17_upstream_read;
  wire    [ 31: 0] std_2s60_burst_17_upstream_readdata_from_sa;
  wire             std_2s60_burst_17_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_17_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_17_upstream_selected_burstcount;
  reg              std_2s60_burst_17_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_17_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_17_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_17_upstream_transaction_burst_count;
  wire             std_2s60_burst_17_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_17_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_17_upstream_waits_for_read;
  wire             std_2s60_burst_17_upstream_waits_for_write;
  wire             std_2s60_burst_17_upstream_write;
  wire    [ 31: 0] std_2s60_burst_17_upstream_writedata;
  wire             wait_for_std_2s60_burst_17_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_17_upstream_end_xfer;
    end


  assign std_2s60_burst_17_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_17_upstream));
  //assign std_2s60_burst_17_upstream_readdatavalid_from_sa = std_2s60_burst_17_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_17_upstream_readdatavalid_from_sa = std_2s60_burst_17_upstream_readdatavalid;

  //assign std_2s60_burst_17_upstream_readdata_from_sa = std_2s60_burst_17_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_17_upstream_readdata_from_sa = std_2s60_burst_17_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_17_upstream = ({cpu_data_master_address_to_slave[25 : 14] , 14'b0} == 26'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_17_upstream_waitrequest_from_sa = std_2s60_burst_17_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_17_upstream_waitrequest_from_sa = std_2s60_burst_17_upstream_waitrequest;

  //std_2s60_burst_17_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_17_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_17_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_17_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_17_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_17_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_17_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_17_upstream;

  //std_2s60_burst_17_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_17_upstream_arb_share_counter_next_value = std_2s60_burst_17_upstream_firsttransfer ? (std_2s60_burst_17_upstream_arb_share_set_values - 1) : |std_2s60_burst_17_upstream_arb_share_counter ? (std_2s60_burst_17_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_17_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_17_upstream_allgrants = |std_2s60_burst_17_upstream_grant_vector;

  //std_2s60_burst_17_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_17_upstream_end_xfer = ~(std_2s60_burst_17_upstream_waits_for_read | std_2s60_burst_17_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream = std_2s60_burst_17_upstream_end_xfer & (~std_2s60_burst_17_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_17_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_17_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream & std_2s60_burst_17_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream & ~std_2s60_burst_17_upstream_non_bursting_master_requests);

  //std_2s60_burst_17_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_17_upstream_arb_counter_enable)
          std_2s60_burst_17_upstream_arb_share_counter <= std_2s60_burst_17_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_17_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_17_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_17_upstream & ~std_2s60_burst_17_upstream_non_bursting_master_requests))
          std_2s60_burst_17_upstream_slavearbiterlockenable <= |std_2s60_burst_17_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_17/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_17_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_17_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_17_upstream_slavearbiterlockenable2 = |std_2s60_burst_17_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_17/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_17_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_17_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_17_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_17_upstream = cpu_data_master_requests_std_2s60_burst_17_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_17_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_17_upstream_move_on_to_next_transaction = std_2s60_burst_17_upstream_this_cycle_is_the_last_burst & std_2s60_burst_17_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_17_upstream, which is an e_mux
  assign std_2s60_burst_17_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_17_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_17_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_17_upstream_module burstcount_fifo_for_std_2s60_burst_17_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_17_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_17_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_17_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_17_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read & std_2s60_burst_17_upstream_load_fifo & ~(std_2s60_burst_17_upstream_this_cycle_is_the_last_burst & std_2s60_burst_17_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_17_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_17_upstream_current_burst_minus_one = std_2s60_burst_17_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_17_upstream, which is an e_mux
  assign std_2s60_burst_17_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read) & ~std_2s60_burst_17_upstream_load_fifo))? std_2s60_burst_17_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read & std_2s60_burst_17_upstream_this_cycle_is_the_last_burst & std_2s60_burst_17_upstream_burstcount_fifo_empty))? std_2s60_burst_17_upstream_selected_burstcount :
    (std_2s60_burst_17_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_17_upstream_transaction_burst_count :
    std_2s60_burst_17_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_17_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_current_burst <= 0;
      else if (std_2s60_burst_17_upstream_readdatavalid_from_sa | (~std_2s60_burst_17_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read)))
          std_2s60_burst_17_upstream_current_burst <= std_2s60_burst_17_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_17_upstream_load_fifo = (~std_2s60_burst_17_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read) & std_2s60_burst_17_upstream_load_fifo))? 1 :
    ~std_2s60_burst_17_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read) & ~std_2s60_burst_17_upstream_load_fifo | std_2s60_burst_17_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_17_upstream_load_fifo <= p0_std_2s60_burst_17_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_17_upstream, which is an e_assign
  assign std_2s60_burst_17_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_17_upstream_current_burst_minus_one) & std_2s60_burst_17_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_17_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_17_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_17_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_17_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_17_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_17_upstream),
      .full                 (),
      .read                 (std_2s60_burst_17_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_17_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_17_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_17_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_17_upstream = std_2s60_burst_17_upstream_readdatavalid_from_sa;

  //std_2s60_burst_17_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_17_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_17/upstream, which is an e_mux
  assign std_2s60_burst_17_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_17_upstream = cpu_data_master_qualified_request_std_2s60_burst_17_upstream;

  //cpu/data_master saved-grant std_2s60_burst_17/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_17_upstream = cpu_data_master_requests_std_2s60_burst_17_upstream;

  //allow new arb cycle for std_2s60_burst_17/upstream, which is an e_assign
  assign std_2s60_burst_17_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_17_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_17_upstream_master_qreq_vector = 1;

  //std_2s60_burst_17_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_17_upstream_firsttransfer = std_2s60_burst_17_upstream_begins_xfer ? std_2s60_burst_17_upstream_unreg_firsttransfer : std_2s60_burst_17_upstream_reg_firsttransfer;

  //std_2s60_burst_17_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_17_upstream_unreg_firsttransfer = ~(std_2s60_burst_17_upstream_slavearbiterlockenable & std_2s60_burst_17_upstream_any_continuerequest);

  //std_2s60_burst_17_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_17_upstream_begins_xfer)
          std_2s60_burst_17_upstream_reg_firsttransfer <= std_2s60_burst_17_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_17_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_17_upstream_next_bbt_burstcount = ((((std_2s60_burst_17_upstream_write) && (std_2s60_burst_17_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_17_upstream_burstcount - 1) :
    ((((std_2s60_burst_17_upstream_read) && (std_2s60_burst_17_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_17_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_17_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_17_upstream_begins_xfer)
          std_2s60_burst_17_upstream_bbt_burstcounter <= std_2s60_burst_17_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_17_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_17_upstream_beginbursttransfer_internal = std_2s60_burst_17_upstream_begins_xfer & (std_2s60_burst_17_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_17_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_17_upstream_read = cpu_data_master_granted_std_2s60_burst_17_upstream & cpu_data_master_read;

  //std_2s60_burst_17_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_17_upstream_write = cpu_data_master_granted_std_2s60_burst_17_upstream & cpu_data_master_write;

  //std_2s60_burst_17_upstream_address mux, which is an e_mux
  assign std_2s60_burst_17_upstream_address = cpu_data_master_address_to_slave;

  //d1_std_2s60_burst_17_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_17_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_17_upstream_end_xfer <= std_2s60_burst_17_upstream_end_xfer;
    end


  //std_2s60_burst_17_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_17_upstream_waits_for_read = std_2s60_burst_17_upstream_in_a_read_cycle & std_2s60_burst_17_upstream_waitrequest_from_sa;

  //std_2s60_burst_17_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_17_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_17_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_17_upstream_in_a_read_cycle;

  //std_2s60_burst_17_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_17_upstream_waits_for_write = std_2s60_burst_17_upstream_in_a_write_cycle & std_2s60_burst_17_upstream_waitrequest_from_sa;

  //std_2s60_burst_17_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_17_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_17_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_17_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_17_upstream_counter = 0;
  //std_2s60_burst_17_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_17_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_17_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_17_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_17_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_17_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_17_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_17/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_17_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_17/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_17_downstream_arbitrator (
                                                 // inputs:
                                                  ad_buf_s1_readdata_from_sa,
                                                  ad_buf_s1_waitrequest_from_sa,
                                                  clk,
                                                  d1_ad_buf_s1_end_xfer,
                                                  reset_n,
                                                  std_2s60_burst_17_downstream_address,
                                                  std_2s60_burst_17_downstream_burstcount,
                                                  std_2s60_burst_17_downstream_byteenable,
                                                  std_2s60_burst_17_downstream_granted_ad_buf_s1,
                                                  std_2s60_burst_17_downstream_qualified_request_ad_buf_s1,
                                                  std_2s60_burst_17_downstream_read,
                                                  std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1,
                                                  std_2s60_burst_17_downstream_requests_ad_buf_s1,
                                                  std_2s60_burst_17_downstream_write,
                                                  std_2s60_burst_17_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_17_downstream_address_to_slave,
                                                  std_2s60_burst_17_downstream_latency_counter,
                                                  std_2s60_burst_17_downstream_readdata,
                                                  std_2s60_burst_17_downstream_readdatavalid,
                                                  std_2s60_burst_17_downstream_reset_n,
                                                  std_2s60_burst_17_downstream_waitrequest
                                               )
;

  output  [ 13: 0] std_2s60_burst_17_downstream_address_to_slave;
  output           std_2s60_burst_17_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_17_downstream_readdata;
  output           std_2s60_burst_17_downstream_readdatavalid;
  output           std_2s60_burst_17_downstream_reset_n;
  output           std_2s60_burst_17_downstream_waitrequest;
  input   [ 31: 0] ad_buf_s1_readdata_from_sa;
  input            ad_buf_s1_waitrequest_from_sa;
  input            clk;
  input            d1_ad_buf_s1_end_xfer;
  input            reset_n;
  input   [ 13: 0] std_2s60_burst_17_downstream_address;
  input            std_2s60_burst_17_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_17_downstream_byteenable;
  input            std_2s60_burst_17_downstream_granted_ad_buf_s1;
  input            std_2s60_burst_17_downstream_qualified_request_ad_buf_s1;
  input            std_2s60_burst_17_downstream_read;
  input            std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1;
  input            std_2s60_burst_17_downstream_requests_ad_buf_s1;
  input            std_2s60_burst_17_downstream_write;
  input   [ 31: 0] std_2s60_burst_17_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_17_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_17_downstream_readdatavalid;
  wire             r_0;
  reg     [ 13: 0] std_2s60_burst_17_downstream_address_last_time;
  wire    [ 13: 0] std_2s60_burst_17_downstream_address_to_slave;
  reg              std_2s60_burst_17_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_17_downstream_byteenable_last_time;
  wire             std_2s60_burst_17_downstream_is_granted_some_slave;
  reg              std_2s60_burst_17_downstream_latency_counter;
  reg              std_2s60_burst_17_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_17_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_17_downstream_readdata;
  wire             std_2s60_burst_17_downstream_readdatavalid;
  wire             std_2s60_burst_17_downstream_reset_n;
  wire             std_2s60_burst_17_downstream_run;
  wire             std_2s60_burst_17_downstream_waitrequest;
  reg              std_2s60_burst_17_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_17_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 | ~std_2s60_burst_17_downstream_requests_ad_buf_s1) & (std_2s60_burst_17_downstream_granted_ad_buf_s1 | ~std_2s60_burst_17_downstream_qualified_request_ad_buf_s1) & ((~std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 | ~(std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write) | (1 & ~ad_buf_s1_waitrequest_from_sa & (std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write)))) & ((~std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 | ~(std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write) | (1 & ~ad_buf_s1_waitrequest_from_sa & (std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_17_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_17_downstream_address_to_slave = std_2s60_burst_17_downstream_address;

  //std_2s60_burst_17_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_17_downstream_read_but_no_slave_selected <= std_2s60_burst_17_downstream_read & std_2s60_burst_17_downstream_run & ~std_2s60_burst_17_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_17_downstream_is_granted_some_slave = std_2s60_burst_17_downstream_granted_ad_buf_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_17_downstream_readdatavalid = std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_17_downstream_readdatavalid = std_2s60_burst_17_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_17_downstream_readdatavalid;

  //std_2s60_burst_17/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_17_downstream_readdata = ad_buf_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_17_downstream_waitrequest = ~std_2s60_burst_17_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_17_downstream_latency_counter <= p1_std_2s60_burst_17_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_17_downstream_latency_counter = ((std_2s60_burst_17_downstream_run & std_2s60_burst_17_downstream_read))? latency_load_value :
    (std_2s60_burst_17_downstream_latency_counter)? std_2s60_burst_17_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {std_2s60_burst_17_downstream_requests_ad_buf_s1}} & 1;

  //std_2s60_burst_17_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_17_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_17_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_address_last_time <= std_2s60_burst_17_downstream_address;
    end


  //std_2s60_burst_17/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_17_downstream_waitrequest & (std_2s60_burst_17_downstream_read | std_2s60_burst_17_downstream_write);
    end


  //std_2s60_burst_17_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_address != std_2s60_burst_17_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_17_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_burstcount_last_time <= std_2s60_burst_17_downstream_burstcount;
    end


  //std_2s60_burst_17_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_burstcount != std_2s60_burst_17_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_17_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_byteenable_last_time <= std_2s60_burst_17_downstream_byteenable;
    end


  //std_2s60_burst_17_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_byteenable != std_2s60_burst_17_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_17_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_read_last_time <= std_2s60_burst_17_downstream_read;
    end


  //std_2s60_burst_17_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_read != std_2s60_burst_17_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_17_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_write_last_time <= std_2s60_burst_17_downstream_write;
    end


  //std_2s60_burst_17_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_write != std_2s60_burst_17_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_17_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_17_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_17_downstream_writedata_last_time <= std_2s60_burst_17_downstream_writedata;
    end


  //std_2s60_burst_17_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_17_downstream_writedata != std_2s60_burst_17_downstream_writedata_last_time) & std_2s60_burst_17_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_17_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_18_upstream_module (
                                                               // inputs:
                                                                clear_fifo,
                                                                clk,
                                                                data_in,
                                                                read,
                                                                reset_n,
                                                                sync_reset,
                                                                write,

                                                               // outputs:
                                                                data_out,
                                                                empty,
                                                                fifo_contains_ones_n,
                                                                full
                                                             )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_18_upstream_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_18_upstream_arbitrator (
                                               // inputs:
                                                clk,
                                                cpu_instruction_master_address_to_slave,
                                                cpu_instruction_master_burstcount,
                                                cpu_instruction_master_latency_counter,
                                                cpu_instruction_master_read,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                                reset_n,
                                                std_2s60_burst_18_upstream_readdata,
                                                std_2s60_burst_18_upstream_readdatavalid,
                                                std_2s60_burst_18_upstream_waitrequest,

                                               // outputs:
                                                cpu_instruction_master_granted_std_2s60_burst_18_upstream,
                                                cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream,
                                                cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                                cpu_instruction_master_requests_std_2s60_burst_18_upstream,
                                                d1_std_2s60_burst_18_upstream_end_xfer,
                                                std_2s60_burst_18_upstream_address,
                                                std_2s60_burst_18_upstream_byteaddress,
                                                std_2s60_burst_18_upstream_byteenable,
                                                std_2s60_burst_18_upstream_debugaccess,
                                                std_2s60_burst_18_upstream_read,
                                                std_2s60_burst_18_upstream_readdata_from_sa,
                                                std_2s60_burst_18_upstream_waitrequest_from_sa,
                                                std_2s60_burst_18_upstream_write
                                             )
;

  output           cpu_instruction_master_granted_std_2s60_burst_18_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_18_upstream;
  output           d1_std_2s60_burst_18_upstream_end_xfer;
  output  [ 13: 0] std_2s60_burst_18_upstream_address;
  output  [ 15: 0] std_2s60_burst_18_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_18_upstream_byteenable;
  output           std_2s60_burst_18_upstream_debugaccess;
  output           std_2s60_burst_18_upstream_read;
  output  [ 31: 0] std_2s60_burst_18_upstream_readdata_from_sa;
  output           std_2s60_burst_18_upstream_waitrequest_from_sa;
  output           std_2s60_burst_18_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_18_upstream_readdata;
  input            std_2s60_burst_18_upstream_readdatavalid;
  input            std_2s60_burst_18_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_18_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_18_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_18_upstream_load_fifo;
  wire    [ 13: 0] std_2s60_burst_18_upstream_address;
  wire             std_2s60_burst_18_upstream_allgrants;
  wire             std_2s60_burst_18_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_18_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_18_upstream_any_continuerequest;
  wire             std_2s60_burst_18_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_18_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_18_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_18_upstream_arb_share_set_values;
  wire             std_2s60_burst_18_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_18_upstream_begins_xfer;
  wire             std_2s60_burst_18_upstream_burstcount_fifo_empty;
  wire    [ 15: 0] std_2s60_burst_18_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_18_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_18_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_18_upstream_current_burst_minus_one;
  wire             std_2s60_burst_18_upstream_debugaccess;
  wire             std_2s60_burst_18_upstream_end_xfer;
  wire             std_2s60_burst_18_upstream_firsttransfer;
  wire             std_2s60_burst_18_upstream_grant_vector;
  wire             std_2s60_burst_18_upstream_in_a_read_cycle;
  wire             std_2s60_burst_18_upstream_in_a_write_cycle;
  reg              std_2s60_burst_18_upstream_load_fifo;
  wire             std_2s60_burst_18_upstream_master_qreq_vector;
  wire             std_2s60_burst_18_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_18_upstream_next_burst_count;
  wire             std_2s60_burst_18_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_18_upstream_read;
  wire    [ 31: 0] std_2s60_burst_18_upstream_readdata_from_sa;
  wire             std_2s60_burst_18_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_18_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_18_upstream_selected_burstcount;
  reg              std_2s60_burst_18_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_18_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_18_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_18_upstream_transaction_burst_count;
  wire             std_2s60_burst_18_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_18_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_18_upstream_waits_for_read;
  wire             std_2s60_burst_18_upstream_waits_for_write;
  wire             std_2s60_burst_18_upstream_write;
  wire             wait_for_std_2s60_burst_18_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_18_upstream_end_xfer;
    end


  assign std_2s60_burst_18_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream));
  //assign std_2s60_burst_18_upstream_readdatavalid_from_sa = std_2s60_burst_18_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_18_upstream_readdatavalid_from_sa = std_2s60_burst_18_upstream_readdatavalid;

  //assign std_2s60_burst_18_upstream_readdata_from_sa = std_2s60_burst_18_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_18_upstream_readdata_from_sa = std_2s60_burst_18_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_18_upstream = (({cpu_instruction_master_address_to_slave[25 : 14] , 14'b0} == 26'h0) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_18_upstream_waitrequest_from_sa = std_2s60_burst_18_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_18_upstream_waitrequest_from_sa = std_2s60_burst_18_upstream_waitrequest;

  //std_2s60_burst_18_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_18_upstream_arb_share_set_values = 1;

  //std_2s60_burst_18_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_18_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_18_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_18_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_18_upstream;

  //std_2s60_burst_18_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_18_upstream_arb_share_counter_next_value = std_2s60_burst_18_upstream_firsttransfer ? (std_2s60_burst_18_upstream_arb_share_set_values - 1) : |std_2s60_burst_18_upstream_arb_share_counter ? (std_2s60_burst_18_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_18_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_18_upstream_allgrants = |std_2s60_burst_18_upstream_grant_vector;

  //std_2s60_burst_18_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_18_upstream_end_xfer = ~(std_2s60_burst_18_upstream_waits_for_read | std_2s60_burst_18_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream = std_2s60_burst_18_upstream_end_xfer & (~std_2s60_burst_18_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_18_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_18_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream & std_2s60_burst_18_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream & ~std_2s60_burst_18_upstream_non_bursting_master_requests);

  //std_2s60_burst_18_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_18_upstream_arb_counter_enable)
          std_2s60_burst_18_upstream_arb_share_counter <= std_2s60_burst_18_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_18_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_18_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_18_upstream & ~std_2s60_burst_18_upstream_non_bursting_master_requests))
          std_2s60_burst_18_upstream_slavearbiterlockenable <= |std_2s60_burst_18_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_18/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_18_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_18_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_18_upstream_slavearbiterlockenable2 = |std_2s60_burst_18_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_18/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_18_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_18_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_18_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream = cpu_instruction_master_requests_std_2s60_burst_18_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_18_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_18_upstream_move_on_to_next_transaction = std_2s60_burst_18_upstream_this_cycle_is_the_last_burst & std_2s60_burst_18_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_18_upstream, which is an e_mux
  assign std_2s60_burst_18_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_18_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_18_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_18_upstream_module burstcount_fifo_for_std_2s60_burst_18_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_18_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_18_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_18_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_18_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read & std_2s60_burst_18_upstream_load_fifo & ~(std_2s60_burst_18_upstream_this_cycle_is_the_last_burst & std_2s60_burst_18_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_18_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_18_upstream_current_burst_minus_one = std_2s60_burst_18_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_18_upstream, which is an e_mux
  assign std_2s60_burst_18_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read) & ~std_2s60_burst_18_upstream_load_fifo))? std_2s60_burst_18_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read & std_2s60_burst_18_upstream_this_cycle_is_the_last_burst & std_2s60_burst_18_upstream_burstcount_fifo_empty))? std_2s60_burst_18_upstream_selected_burstcount :
    (std_2s60_burst_18_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_18_upstream_transaction_burst_count :
    std_2s60_burst_18_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_18_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_upstream_current_burst <= 0;
      else if (std_2s60_burst_18_upstream_readdatavalid_from_sa | (~std_2s60_burst_18_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read)))
          std_2s60_burst_18_upstream_current_burst <= std_2s60_burst_18_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_18_upstream_load_fifo = (~std_2s60_burst_18_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read) & std_2s60_burst_18_upstream_load_fifo))? 1 :
    ~std_2s60_burst_18_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read) & ~std_2s60_burst_18_upstream_load_fifo | std_2s60_burst_18_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_18_upstream_load_fifo <= p0_std_2s60_burst_18_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_18_upstream, which is an e_assign
  assign std_2s60_burst_18_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_18_upstream_current_burst_minus_one) & std_2s60_burst_18_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_18_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_18_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_18_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_18_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_18_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_18_upstream),
      .full                 (),
      .read                 (std_2s60_burst_18_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_18_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_18_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream = std_2s60_burst_18_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_18/upstream, which is an e_mux
  assign std_2s60_burst_18_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_18_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_18/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_18_upstream = cpu_instruction_master_requests_std_2s60_burst_18_upstream;

  //allow new arb cycle for std_2s60_burst_18/upstream, which is an e_assign
  assign std_2s60_burst_18_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_18_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_18_upstream_master_qreq_vector = 1;

  //std_2s60_burst_18_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_18_upstream_firsttransfer = std_2s60_burst_18_upstream_begins_xfer ? std_2s60_burst_18_upstream_unreg_firsttransfer : std_2s60_burst_18_upstream_reg_firsttransfer;

  //std_2s60_burst_18_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_18_upstream_unreg_firsttransfer = ~(std_2s60_burst_18_upstream_slavearbiterlockenable & std_2s60_burst_18_upstream_any_continuerequest);

  //std_2s60_burst_18_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_18_upstream_begins_xfer)
          std_2s60_burst_18_upstream_reg_firsttransfer <= std_2s60_burst_18_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_18_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_18_upstream_beginbursttransfer_internal = std_2s60_burst_18_upstream_begins_xfer;

  //std_2s60_burst_18_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_18_upstream_read = cpu_instruction_master_granted_std_2s60_burst_18_upstream & cpu_instruction_master_read;

  //std_2s60_burst_18_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_18_upstream_write = 0;

  //std_2s60_burst_18_upstream_address mux, which is an e_mux
  assign std_2s60_burst_18_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_std_2s60_burst_18_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_18_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_18_upstream_end_xfer <= std_2s60_burst_18_upstream_end_xfer;
    end


  //std_2s60_burst_18_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_18_upstream_waits_for_read = std_2s60_burst_18_upstream_in_a_read_cycle & std_2s60_burst_18_upstream_waitrequest_from_sa;

  //std_2s60_burst_18_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_18_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_18_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_18_upstream_in_a_read_cycle;

  //std_2s60_burst_18_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_18_upstream_waits_for_write = std_2s60_burst_18_upstream_in_a_write_cycle & std_2s60_burst_18_upstream_waitrequest_from_sa;

  //std_2s60_burst_18_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_18_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_18_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_18_upstream_counter = 0;
  //std_2s60_burst_18_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_18_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_18_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_18/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_18_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_18/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_18_downstream_arbitrator (
                                                 // inputs:
                                                  ad_buf_s1_readdata_from_sa,
                                                  ad_buf_s1_waitrequest_from_sa,
                                                  clk,
                                                  d1_ad_buf_s1_end_xfer,
                                                  reset_n,
                                                  std_2s60_burst_18_downstream_address,
                                                  std_2s60_burst_18_downstream_burstcount,
                                                  std_2s60_burst_18_downstream_byteenable,
                                                  std_2s60_burst_18_downstream_granted_ad_buf_s1,
                                                  std_2s60_burst_18_downstream_qualified_request_ad_buf_s1,
                                                  std_2s60_burst_18_downstream_read,
                                                  std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1,
                                                  std_2s60_burst_18_downstream_requests_ad_buf_s1,
                                                  std_2s60_burst_18_downstream_write,
                                                  std_2s60_burst_18_downstream_writedata,

                                                 // outputs:
                                                  std_2s60_burst_18_downstream_address_to_slave,
                                                  std_2s60_burst_18_downstream_latency_counter,
                                                  std_2s60_burst_18_downstream_readdata,
                                                  std_2s60_burst_18_downstream_readdatavalid,
                                                  std_2s60_burst_18_downstream_reset_n,
                                                  std_2s60_burst_18_downstream_waitrequest
                                               )
;

  output  [ 13: 0] std_2s60_burst_18_downstream_address_to_slave;
  output           std_2s60_burst_18_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_18_downstream_readdata;
  output           std_2s60_burst_18_downstream_readdatavalid;
  output           std_2s60_burst_18_downstream_reset_n;
  output           std_2s60_burst_18_downstream_waitrequest;
  input   [ 31: 0] ad_buf_s1_readdata_from_sa;
  input            ad_buf_s1_waitrequest_from_sa;
  input            clk;
  input            d1_ad_buf_s1_end_xfer;
  input            reset_n;
  input   [ 13: 0] std_2s60_burst_18_downstream_address;
  input            std_2s60_burst_18_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_18_downstream_byteenable;
  input            std_2s60_burst_18_downstream_granted_ad_buf_s1;
  input            std_2s60_burst_18_downstream_qualified_request_ad_buf_s1;
  input            std_2s60_burst_18_downstream_read;
  input            std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1;
  input            std_2s60_burst_18_downstream_requests_ad_buf_s1;
  input            std_2s60_burst_18_downstream_write;
  input   [ 31: 0] std_2s60_burst_18_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_18_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_18_downstream_readdatavalid;
  wire             r_0;
  reg     [ 13: 0] std_2s60_burst_18_downstream_address_last_time;
  wire    [ 13: 0] std_2s60_burst_18_downstream_address_to_slave;
  reg              std_2s60_burst_18_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_18_downstream_byteenable_last_time;
  wire             std_2s60_burst_18_downstream_is_granted_some_slave;
  reg              std_2s60_burst_18_downstream_latency_counter;
  reg              std_2s60_burst_18_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_18_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_18_downstream_readdata;
  wire             std_2s60_burst_18_downstream_readdatavalid;
  wire             std_2s60_burst_18_downstream_reset_n;
  wire             std_2s60_burst_18_downstream_run;
  wire             std_2s60_burst_18_downstream_waitrequest;
  reg              std_2s60_burst_18_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_18_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 | ~std_2s60_burst_18_downstream_requests_ad_buf_s1) & (std_2s60_burst_18_downstream_granted_ad_buf_s1 | ~std_2s60_burst_18_downstream_qualified_request_ad_buf_s1) & ((~std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 | ~(std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write) | (1 & ~ad_buf_s1_waitrequest_from_sa & (std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write)))) & ((~std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 | ~(std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write) | (1 & ~ad_buf_s1_waitrequest_from_sa & (std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_18_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_18_downstream_address_to_slave = std_2s60_burst_18_downstream_address;

  //std_2s60_burst_18_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_18_downstream_read_but_no_slave_selected <= std_2s60_burst_18_downstream_read & std_2s60_burst_18_downstream_run & ~std_2s60_burst_18_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_18_downstream_is_granted_some_slave = std_2s60_burst_18_downstream_granted_ad_buf_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_18_downstream_readdatavalid = std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_18_downstream_readdatavalid = std_2s60_burst_18_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_18_downstream_readdatavalid;

  //std_2s60_burst_18/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_18_downstream_readdata = ad_buf_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_18_downstream_waitrequest = ~std_2s60_burst_18_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_18_downstream_latency_counter <= p1_std_2s60_burst_18_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_18_downstream_latency_counter = ((std_2s60_burst_18_downstream_run & std_2s60_burst_18_downstream_read))? latency_load_value :
    (std_2s60_burst_18_downstream_latency_counter)? std_2s60_burst_18_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {std_2s60_burst_18_downstream_requests_ad_buf_s1}} & 1;

  //std_2s60_burst_18_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_18_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_18_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_address_last_time <= std_2s60_burst_18_downstream_address;
    end


  //std_2s60_burst_18/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_18_downstream_waitrequest & (std_2s60_burst_18_downstream_read | std_2s60_burst_18_downstream_write);
    end


  //std_2s60_burst_18_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_address != std_2s60_burst_18_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_18_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_burstcount_last_time <= std_2s60_burst_18_downstream_burstcount;
    end


  //std_2s60_burst_18_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_burstcount != std_2s60_burst_18_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_18_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_byteenable_last_time <= std_2s60_burst_18_downstream_byteenable;
    end


  //std_2s60_burst_18_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_byteenable != std_2s60_burst_18_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_18_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_read_last_time <= std_2s60_burst_18_downstream_read;
    end


  //std_2s60_burst_18_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_read != std_2s60_burst_18_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_18_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_write_last_time <= std_2s60_burst_18_downstream_write;
    end


  //std_2s60_burst_18_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_write != std_2s60_burst_18_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_18_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_18_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_18_downstream_writedata_last_time <= std_2s60_burst_18_downstream_writedata;
    end


  //std_2s60_burst_18_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_18_downstream_writedata != std_2s60_burst_18_downstream_writedata_last_time) & std_2s60_burst_18_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_18_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_2_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  5: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  5: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  5: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  5: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  5: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  5: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  5: 0] p3_stage_3;
  reg     [  5: 0] stage_0;
  reg     [  5: 0] stage_1;
  reg     [  5: 0] stage_2;
  reg     [  5: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_2_upstream_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_2_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_instruction_master_address_to_slave,
                                               cpu_instruction_master_burstcount,
                                               cpu_instruction_master_dbs_address,
                                               cpu_instruction_master_latency_counter,
                                               cpu_instruction_master_read,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                               reset_n,
                                               std_2s60_burst_2_upstream_readdata,
                                               std_2s60_burst_2_upstream_readdatavalid,
                                               std_2s60_burst_2_upstream_waitrequest,

                                              // outputs:
                                               cpu_instruction_master_granted_std_2s60_burst_2_upstream,
                                               cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                               cpu_instruction_master_requests_std_2s60_burst_2_upstream,
                                               d1_std_2s60_burst_2_upstream_end_xfer,
                                               std_2s60_burst_2_upstream_address,
                                               std_2s60_burst_2_upstream_byteaddress,
                                               std_2s60_burst_2_upstream_byteenable,
                                               std_2s60_burst_2_upstream_debugaccess,
                                               std_2s60_burst_2_upstream_read,
                                               std_2s60_burst_2_upstream_readdata_from_sa,
                                               std_2s60_burst_2_upstream_waitrequest_from_sa,
                                               std_2s60_burst_2_upstream_write
                                            )
;

  output           cpu_instruction_master_granted_std_2s60_burst_2_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_2_upstream;
  output           d1_std_2s60_burst_2_upstream_end_xfer;
  output  [ 23: 0] std_2s60_burst_2_upstream_address;
  output  [ 23: 0] std_2s60_burst_2_upstream_byteaddress;
  output           std_2s60_burst_2_upstream_byteenable;
  output           std_2s60_burst_2_upstream_debugaccess;
  output           std_2s60_burst_2_upstream_read;
  output  [  7: 0] std_2s60_burst_2_upstream_readdata_from_sa;
  output           std_2s60_burst_2_upstream_waitrequest_from_sa;
  output           std_2s60_burst_2_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input   [  1: 0] cpu_instruction_master_dbs_address;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [  7: 0] std_2s60_burst_2_upstream_readdata;
  input            std_2s60_burst_2_upstream_readdatavalid;
  input            std_2s60_burst_2_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_2_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_2_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_2_upstream_load_fifo;
  wire    [ 23: 0] std_2s60_burst_2_upstream_address;
  wire             std_2s60_burst_2_upstream_allgrants;
  wire             std_2s60_burst_2_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_2_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_2_upstream_any_continuerequest;
  wire             std_2s60_burst_2_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_2_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_2_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_2_upstream_arb_share_set_values;
  wire             std_2s60_burst_2_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_2_upstream_begins_xfer;
  wire             std_2s60_burst_2_upstream_burstcount_fifo_empty;
  wire    [ 23: 0] std_2s60_burst_2_upstream_byteaddress;
  wire             std_2s60_burst_2_upstream_byteenable;
  reg     [  5: 0] std_2s60_burst_2_upstream_current_burst;
  wire    [  5: 0] std_2s60_burst_2_upstream_current_burst_minus_one;
  wire             std_2s60_burst_2_upstream_debugaccess;
  wire             std_2s60_burst_2_upstream_end_xfer;
  wire             std_2s60_burst_2_upstream_firsttransfer;
  wire             std_2s60_burst_2_upstream_grant_vector;
  wire             std_2s60_burst_2_upstream_in_a_read_cycle;
  wire             std_2s60_burst_2_upstream_in_a_write_cycle;
  reg              std_2s60_burst_2_upstream_load_fifo;
  wire             std_2s60_burst_2_upstream_master_qreq_vector;
  wire             std_2s60_burst_2_upstream_move_on_to_next_transaction;
  wire    [  5: 0] std_2s60_burst_2_upstream_next_burst_count;
  wire             std_2s60_burst_2_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_2_upstream_read;
  wire    [  7: 0] std_2s60_burst_2_upstream_readdata_from_sa;
  wire             std_2s60_burst_2_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_2_upstream_reg_firsttransfer;
  wire    [  5: 0] std_2s60_burst_2_upstream_selected_burstcount;
  reg              std_2s60_burst_2_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_2_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_2_upstream_this_cycle_is_the_last_burst;
  wire    [  5: 0] std_2s60_burst_2_upstream_transaction_burst_count;
  wire             std_2s60_burst_2_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_2_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_2_upstream_waits_for_read;
  wire             std_2s60_burst_2_upstream_waits_for_write;
  wire             std_2s60_burst_2_upstream_write;
  wire             wait_for_std_2s60_burst_2_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_2_upstream_end_xfer;
    end


  assign std_2s60_burst_2_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream));
  //assign std_2s60_burst_2_upstream_readdatavalid_from_sa = std_2s60_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_2_upstream_readdatavalid_from_sa = std_2s60_burst_2_upstream_readdatavalid;

  //assign std_2s60_burst_2_upstream_readdata_from_sa = std_2s60_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_2_upstream_readdata_from_sa = std_2s60_burst_2_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_2_upstream = (({cpu_instruction_master_address_to_slave[25 : 24] , 24'b0} == 26'h3000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_2_upstream_waitrequest_from_sa = std_2s60_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_2_upstream_waitrequest_from_sa = std_2s60_burst_2_upstream_waitrequest;

  //std_2s60_burst_2_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_2_upstream_arb_share_set_values = 1;

  //std_2s60_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_2_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_2_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_2_upstream;

  //std_2s60_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_2_upstream_arb_share_counter_next_value = std_2s60_burst_2_upstream_firsttransfer ? (std_2s60_burst_2_upstream_arb_share_set_values - 1) : |std_2s60_burst_2_upstream_arb_share_counter ? (std_2s60_burst_2_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_2_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_2_upstream_allgrants = |std_2s60_burst_2_upstream_grant_vector;

  //std_2s60_burst_2_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_2_upstream_end_xfer = ~(std_2s60_burst_2_upstream_waits_for_read | std_2s60_burst_2_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream = std_2s60_burst_2_upstream_end_xfer & (~std_2s60_burst_2_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_2_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream & std_2s60_burst_2_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream & ~std_2s60_burst_2_upstream_non_bursting_master_requests);

  //std_2s60_burst_2_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_2_upstream_arb_counter_enable)
          std_2s60_burst_2_upstream_arb_share_counter <= std_2s60_burst_2_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_2_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_2_upstream & ~std_2s60_burst_2_upstream_non_bursting_master_requests))
          std_2s60_burst_2_upstream_slavearbiterlockenable <= |std_2s60_burst_2_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_2/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_2_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_2_upstream_slavearbiterlockenable2 = |std_2s60_burst_2_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_2/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_2_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_2_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream = cpu_instruction_master_requests_std_2s60_burst_2_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_2_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_2_upstream_move_on_to_next_transaction = std_2s60_burst_2_upstream_this_cycle_is_the_last_burst & std_2s60_burst_2_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_2_upstream, which is an e_mux
  assign std_2s60_burst_2_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_2_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_2_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_2_upstream_module burstcount_fifo_for_std_2s60_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_2_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_2_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_2_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_2_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read & std_2s60_burst_2_upstream_load_fifo & ~(std_2s60_burst_2_upstream_this_cycle_is_the_last_burst & std_2s60_burst_2_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_2_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_2_upstream_current_burst_minus_one = std_2s60_burst_2_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_2_upstream, which is an e_mux
  assign std_2s60_burst_2_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read) & ~std_2s60_burst_2_upstream_load_fifo))? {std_2s60_burst_2_upstream_selected_burstcount, 2'b0} :
    ((in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read & std_2s60_burst_2_upstream_this_cycle_is_the_last_burst & std_2s60_burst_2_upstream_burstcount_fifo_empty))? {std_2s60_burst_2_upstream_selected_burstcount, 2'b0} :
    (std_2s60_burst_2_upstream_this_cycle_is_the_last_burst)? {std_2s60_burst_2_upstream_transaction_burst_count,  2'b0} :
    std_2s60_burst_2_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_2_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_upstream_current_burst <= 0;
      else if (std_2s60_burst_2_upstream_readdatavalid_from_sa | (~std_2s60_burst_2_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read)))
          std_2s60_burst_2_upstream_current_burst <= std_2s60_burst_2_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_2_upstream_load_fifo = (~std_2s60_burst_2_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read) & std_2s60_burst_2_upstream_load_fifo))? 1 :
    ~std_2s60_burst_2_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read) & ~std_2s60_burst_2_upstream_load_fifo | std_2s60_burst_2_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_2_upstream_load_fifo <= p0_std_2s60_burst_2_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_2_upstream, which is an e_assign
  assign std_2s60_burst_2_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_2_upstream_current_burst_minus_one) & std_2s60_burst_2_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_2_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_2_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_2_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_2_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_2_upstream),
      .full                 (),
      .read                 (std_2s60_burst_2_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_2_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_2_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream = std_2s60_burst_2_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_2/upstream, which is an e_mux
  assign std_2s60_burst_2_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_2_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_2/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_2_upstream = cpu_instruction_master_requests_std_2s60_burst_2_upstream;

  //allow new arb cycle for std_2s60_burst_2/upstream, which is an e_assign
  assign std_2s60_burst_2_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_2_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_2_upstream_master_qreq_vector = 1;

  //std_2s60_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_2_upstream_firsttransfer = std_2s60_burst_2_upstream_begins_xfer ? std_2s60_burst_2_upstream_unreg_firsttransfer : std_2s60_burst_2_upstream_reg_firsttransfer;

  //std_2s60_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_2_upstream_unreg_firsttransfer = ~(std_2s60_burst_2_upstream_slavearbiterlockenable & std_2s60_burst_2_upstream_any_continuerequest);

  //std_2s60_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_2_upstream_begins_xfer)
          std_2s60_burst_2_upstream_reg_firsttransfer <= std_2s60_burst_2_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_2_upstream_beginbursttransfer_internal = std_2s60_burst_2_upstream_begins_xfer;

  //std_2s60_burst_2_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_2_upstream_read = cpu_instruction_master_granted_std_2s60_burst_2_upstream & cpu_instruction_master_read;

  //std_2s60_burst_2_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_2_upstream_write = 0;

  //std_2s60_burst_2_upstream_address mux, which is an e_mux
  assign std_2s60_burst_2_upstream_address = {cpu_instruction_master_address_to_slave >> 2,
    cpu_instruction_master_dbs_address[1 : 0]};

  //d1_std_2s60_burst_2_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_2_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_2_upstream_end_xfer <= std_2s60_burst_2_upstream_end_xfer;
    end


  //std_2s60_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_2_upstream_waits_for_read = std_2s60_burst_2_upstream_in_a_read_cycle & std_2s60_burst_2_upstream_waitrequest_from_sa;

  //std_2s60_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_2_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_2_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_2_upstream_in_a_read_cycle;

  //std_2s60_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_2_upstream_waits_for_write = std_2s60_burst_2_upstream_in_a_write_cycle & std_2s60_burst_2_upstream_waitrequest_from_sa;

  //std_2s60_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_2_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_2_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_2_upstream_counter = 0;
  //std_2s60_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_2_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_2_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_2/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_2_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_2/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_2_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_flash_bus_avalon_slave_end_xfer,
                                                 ext_flash_s1_wait_counter_eq_0,
                                                 incoming_ext_flash_bus_data_with_Xs_converted_to_0,
                                                 reset_n,
                                                 std_2s60_burst_2_downstream_address,
                                                 std_2s60_burst_2_downstream_burstcount,
                                                 std_2s60_burst_2_downstream_byteenable,
                                                 std_2s60_burst_2_downstream_granted_ext_flash_s1,
                                                 std_2s60_burst_2_downstream_qualified_request_ext_flash_s1,
                                                 std_2s60_burst_2_downstream_read,
                                                 std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1,
                                                 std_2s60_burst_2_downstream_requests_ext_flash_s1,
                                                 std_2s60_burst_2_downstream_write,
                                                 std_2s60_burst_2_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_2_downstream_address_to_slave,
                                                 std_2s60_burst_2_downstream_latency_counter,
                                                 std_2s60_burst_2_downstream_readdata,
                                                 std_2s60_burst_2_downstream_readdatavalid,
                                                 std_2s60_burst_2_downstream_reset_n,
                                                 std_2s60_burst_2_downstream_waitrequest
                                              )
;

  output  [ 23: 0] std_2s60_burst_2_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_2_downstream_latency_counter;
  output  [  7: 0] std_2s60_burst_2_downstream_readdata;
  output           std_2s60_burst_2_downstream_readdatavalid;
  output           std_2s60_burst_2_downstream_reset_n;
  output           std_2s60_burst_2_downstream_waitrequest;
  input            clk;
  input            d1_ext_flash_bus_avalon_slave_end_xfer;
  input            ext_flash_s1_wait_counter_eq_0;
  input   [  7: 0] incoming_ext_flash_bus_data_with_Xs_converted_to_0;
  input            reset_n;
  input   [ 23: 0] std_2s60_burst_2_downstream_address;
  input            std_2s60_burst_2_downstream_burstcount;
  input            std_2s60_burst_2_downstream_byteenable;
  input            std_2s60_burst_2_downstream_granted_ext_flash_s1;
  input            std_2s60_burst_2_downstream_qualified_request_ext_flash_s1;
  input            std_2s60_burst_2_downstream_read;
  input            std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1;
  input            std_2s60_burst_2_downstream_requests_ext_flash_s1;
  input            std_2s60_burst_2_downstream_write;
  input   [  7: 0] std_2s60_burst_2_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_2_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_2_downstream_readdatavalid;
  wire             r_0;
  reg     [ 23: 0] std_2s60_burst_2_downstream_address_last_time;
  wire    [ 23: 0] std_2s60_burst_2_downstream_address_to_slave;
  reg              std_2s60_burst_2_downstream_burstcount_last_time;
  reg              std_2s60_burst_2_downstream_byteenable_last_time;
  wire             std_2s60_burst_2_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_2_downstream_latency_counter;
  reg              std_2s60_burst_2_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_2_downstream_read_last_time;
  wire    [  7: 0] std_2s60_burst_2_downstream_readdata;
  wire             std_2s60_burst_2_downstream_readdatavalid;
  wire             std_2s60_burst_2_downstream_reset_n;
  wire             std_2s60_burst_2_downstream_run;
  wire             std_2s60_burst_2_downstream_waitrequest;
  reg              std_2s60_burst_2_downstream_write_last_time;
  reg     [  7: 0] std_2s60_burst_2_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_2_downstream_requests_ext_flash_s1) & (std_2s60_burst_2_downstream_granted_ext_flash_s1 | ~std_2s60_burst_2_downstream_qualified_request_ext_flash_s1) & ((~std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_2_downstream_read | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_ext_flash_bus_avalon_slave_end_xfer)) & std_2s60_burst_2_downstream_read))) & ((~std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_2_downstream_write | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_ext_flash_bus_avalon_slave_end_xfer)) & std_2s60_burst_2_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_2_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_2_downstream_address_to_slave = std_2s60_burst_2_downstream_address;

  //std_2s60_burst_2_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_2_downstream_read_but_no_slave_selected <= std_2s60_burst_2_downstream_read & std_2s60_burst_2_downstream_run & ~std_2s60_burst_2_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_2_downstream_is_granted_some_slave = std_2s60_burst_2_downstream_granted_ext_flash_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_2_downstream_readdatavalid = std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_2_downstream_readdatavalid = std_2s60_burst_2_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_2_downstream_readdatavalid;

  //std_2s60_burst_2/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_2_downstream_readdata = incoming_ext_flash_bus_data_with_Xs_converted_to_0;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_2_downstream_waitrequest = ~std_2s60_burst_2_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_2_downstream_latency_counter <= p1_std_2s60_burst_2_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_2_downstream_latency_counter = ((std_2s60_burst_2_downstream_run & std_2s60_burst_2_downstream_read))? latency_load_value :
    (std_2s60_burst_2_downstream_latency_counter)? std_2s60_burst_2_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {2 {std_2s60_burst_2_downstream_requests_ext_flash_s1}} & 2;

  //std_2s60_burst_2_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_2_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_2_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_address_last_time <= std_2s60_burst_2_downstream_address;
    end


  //std_2s60_burst_2/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_2_downstream_waitrequest & (std_2s60_burst_2_downstream_read | std_2s60_burst_2_downstream_write);
    end


  //std_2s60_burst_2_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_address != std_2s60_burst_2_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_2_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_burstcount_last_time <= std_2s60_burst_2_downstream_burstcount;
    end


  //std_2s60_burst_2_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_burstcount != std_2s60_burst_2_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_2_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_byteenable_last_time <= std_2s60_burst_2_downstream_byteenable;
    end


  //std_2s60_burst_2_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_byteenable != std_2s60_burst_2_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_2_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_read_last_time <= std_2s60_burst_2_downstream_read;
    end


  //std_2s60_burst_2_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_read != std_2s60_burst_2_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_2_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_write_last_time <= std_2s60_burst_2_downstream_write;
    end


  //std_2s60_burst_2_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_write != std_2s60_burst_2_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_2_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_2_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_2_downstream_writedata_last_time <= std_2s60_burst_2_downstream_writedata;
    end


  //std_2s60_burst_2_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_2_downstream_writedata != std_2s60_burst_2_downstream_writedata_last_time) & std_2s60_burst_2_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_2_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_3_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  5: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  5: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  5: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  5: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  5: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  5: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  5: 0] p3_stage_3;
  reg     [  5: 0] stage_0;
  reg     [  5: 0] stage_1;
  reg     [  5: 0] stage_2;
  reg     [  5: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_3_upstream_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_3_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_burstcount,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_dbs_address,
                                               cpu_data_master_dbs_write_8,
                                               cpu_data_master_debugaccess,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                               cpu_data_master_write,
                                               reset_n,
                                               std_2s60_burst_3_upstream_readdata,
                                               std_2s60_burst_3_upstream_readdatavalid,
                                               std_2s60_burst_3_upstream_waitrequest,

                                              // outputs:
                                               cpu_data_master_byteenable_std_2s60_burst_3_upstream,
                                               cpu_data_master_granted_std_2s60_burst_3_upstream,
                                               cpu_data_master_qualified_request_std_2s60_burst_3_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                               cpu_data_master_requests_std_2s60_burst_3_upstream,
                                               d1_std_2s60_burst_3_upstream_end_xfer,
                                               std_2s60_burst_3_upstream_address,
                                               std_2s60_burst_3_upstream_burstcount,
                                               std_2s60_burst_3_upstream_byteaddress,
                                               std_2s60_burst_3_upstream_byteenable,
                                               std_2s60_burst_3_upstream_debugaccess,
                                               std_2s60_burst_3_upstream_read,
                                               std_2s60_burst_3_upstream_readdata_from_sa,
                                               std_2s60_burst_3_upstream_waitrequest_from_sa,
                                               std_2s60_burst_3_upstream_write,
                                               std_2s60_burst_3_upstream_writedata
                                            )
;

  output           cpu_data_master_byteenable_std_2s60_burst_3_upstream;
  output           cpu_data_master_granted_std_2s60_burst_3_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_3_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_3_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_3_upstream;
  output           d1_std_2s60_burst_3_upstream_end_xfer;
  output  [ 23: 0] std_2s60_burst_3_upstream_address;
  output  [  3: 0] std_2s60_burst_3_upstream_burstcount;
  output  [ 23: 0] std_2s60_burst_3_upstream_byteaddress;
  output           std_2s60_burst_3_upstream_byteenable;
  output           std_2s60_burst_3_upstream_debugaccess;
  output           std_2s60_burst_3_upstream_read;
  output  [  7: 0] std_2s60_burst_3_upstream_readdata_from_sa;
  output           std_2s60_burst_3_upstream_waitrequest_from_sa;
  output           std_2s60_burst_3_upstream_write;
  output  [  7: 0] std_2s60_burst_3_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_dbs_address;
  input   [  7: 0] cpu_data_master_dbs_write_8;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input            reset_n;
  input   [  7: 0] std_2s60_burst_3_upstream_readdata;
  input            std_2s60_burst_3_upstream_readdatavalid;
  input            std_2s60_burst_3_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_0;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_1;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_2;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_3;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_3_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_3_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_3_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_3_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_3_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_3_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_3_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_3_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_3_upstream_load_fifo;
  wire    [ 23: 0] std_2s60_burst_3_upstream_address;
  wire             std_2s60_burst_3_upstream_allgrants;
  wire             std_2s60_burst_3_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_3_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_3_upstream_any_continuerequest;
  wire             std_2s60_burst_3_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_3_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_3_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_3_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_3_upstream_bbt_burstcounter;
  wire             std_2s60_burst_3_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_3_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_3_upstream_burstcount;
  wire             std_2s60_burst_3_upstream_burstcount_fifo_empty;
  wire    [ 23: 0] std_2s60_burst_3_upstream_byteaddress;
  wire             std_2s60_burst_3_upstream_byteenable;
  reg     [  5: 0] std_2s60_burst_3_upstream_current_burst;
  wire    [  5: 0] std_2s60_burst_3_upstream_current_burst_minus_one;
  wire             std_2s60_burst_3_upstream_debugaccess;
  wire             std_2s60_burst_3_upstream_end_xfer;
  wire             std_2s60_burst_3_upstream_firsttransfer;
  wire             std_2s60_burst_3_upstream_grant_vector;
  wire             std_2s60_burst_3_upstream_in_a_read_cycle;
  wire             std_2s60_burst_3_upstream_in_a_write_cycle;
  reg              std_2s60_burst_3_upstream_load_fifo;
  wire             std_2s60_burst_3_upstream_master_qreq_vector;
  wire             std_2s60_burst_3_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_3_upstream_next_bbt_burstcount;
  wire    [  5: 0] std_2s60_burst_3_upstream_next_burst_count;
  wire             std_2s60_burst_3_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_3_upstream_read;
  wire    [  7: 0] std_2s60_burst_3_upstream_readdata_from_sa;
  wire             std_2s60_burst_3_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_3_upstream_reg_firsttransfer;
  wire    [  5: 0] std_2s60_burst_3_upstream_selected_burstcount;
  reg              std_2s60_burst_3_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_3_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_3_upstream_this_cycle_is_the_last_burst;
  wire    [  5: 0] std_2s60_burst_3_upstream_transaction_burst_count;
  wire             std_2s60_burst_3_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_3_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_3_upstream_waits_for_read;
  wire             std_2s60_burst_3_upstream_waits_for_write;
  wire             std_2s60_burst_3_upstream_write;
  wire    [  7: 0] std_2s60_burst_3_upstream_writedata;
  wire             wait_for_std_2s60_burst_3_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_3_upstream_end_xfer;
    end


  assign std_2s60_burst_3_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_3_upstream));
  //assign std_2s60_burst_3_upstream_readdatavalid_from_sa = std_2s60_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_3_upstream_readdatavalid_from_sa = std_2s60_burst_3_upstream_readdatavalid;

  //assign std_2s60_burst_3_upstream_readdata_from_sa = std_2s60_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_3_upstream_readdata_from_sa = std_2s60_burst_3_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_3_upstream = ({cpu_data_master_address_to_slave[25 : 24] , 24'b0} == 26'h3000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_3_upstream_waitrequest_from_sa = std_2s60_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_3_upstream_waitrequest_from_sa = std_2s60_burst_3_upstream_waitrequest;

  //std_2s60_burst_3_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_3_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_3_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount<< 2 : 1)) :
    1;

  //std_2s60_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_3_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_3_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_3_upstream;

  //std_2s60_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_3_upstream_arb_share_counter_next_value = std_2s60_burst_3_upstream_firsttransfer ? (std_2s60_burst_3_upstream_arb_share_set_values - 1) : |std_2s60_burst_3_upstream_arb_share_counter ? (std_2s60_burst_3_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_3_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_3_upstream_allgrants = |std_2s60_burst_3_upstream_grant_vector;

  //std_2s60_burst_3_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_3_upstream_end_xfer = ~(std_2s60_burst_3_upstream_waits_for_read | std_2s60_burst_3_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream = std_2s60_burst_3_upstream_end_xfer & (~std_2s60_burst_3_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_3_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream & std_2s60_burst_3_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream & ~std_2s60_burst_3_upstream_non_bursting_master_requests);

  //std_2s60_burst_3_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_3_upstream_arb_counter_enable)
          std_2s60_burst_3_upstream_arb_share_counter <= std_2s60_burst_3_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_3_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_3_upstream & ~std_2s60_burst_3_upstream_non_bursting_master_requests))
          std_2s60_burst_3_upstream_slavearbiterlockenable <= |std_2s60_burst_3_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_3/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_3_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_3_upstream_slavearbiterlockenable2 = |std_2s60_burst_3_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_3/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_3_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_3_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_3_upstream = cpu_data_master_requests_std_2s60_burst_3_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_3_upstream_move_on_to_next_transaction = std_2s60_burst_3_upstream_this_cycle_is_the_last_burst & std_2s60_burst_3_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_3_upstream, which is an e_mux
  assign std_2s60_burst_3_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_3_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_3_upstream_module burstcount_fifo_for_std_2s60_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_3_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_3_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_3_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_3_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read & std_2s60_burst_3_upstream_load_fifo & ~(std_2s60_burst_3_upstream_this_cycle_is_the_last_burst & std_2s60_burst_3_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_3_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_3_upstream_current_burst_minus_one = std_2s60_burst_3_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_3_upstream, which is an e_mux
  assign std_2s60_burst_3_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read) & ~std_2s60_burst_3_upstream_load_fifo))? {std_2s60_burst_3_upstream_selected_burstcount, 2'b0} :
    ((in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read & std_2s60_burst_3_upstream_this_cycle_is_the_last_burst & std_2s60_burst_3_upstream_burstcount_fifo_empty))? {std_2s60_burst_3_upstream_selected_burstcount, 2'b0} :
    (std_2s60_burst_3_upstream_this_cycle_is_the_last_burst)? {std_2s60_burst_3_upstream_transaction_burst_count,  2'b0} :
    std_2s60_burst_3_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_3_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_current_burst <= 0;
      else if (std_2s60_burst_3_upstream_readdatavalid_from_sa | (~std_2s60_burst_3_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read)))
          std_2s60_burst_3_upstream_current_burst <= std_2s60_burst_3_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_3_upstream_load_fifo = (~std_2s60_burst_3_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read) & std_2s60_burst_3_upstream_load_fifo))? 1 :
    ~std_2s60_burst_3_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read) & ~std_2s60_burst_3_upstream_load_fifo | std_2s60_burst_3_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_3_upstream_load_fifo <= p0_std_2s60_burst_3_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_3_upstream, which is an e_assign
  assign std_2s60_burst_3_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_3_upstream_current_burst_minus_one) & std_2s60_burst_3_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_3_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_3_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_3_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_3_upstream),
      .full                 (),
      .read                 (std_2s60_burst_3_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_3_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_3_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_3_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_3_upstream = std_2s60_burst_3_upstream_readdatavalid_from_sa;

  //std_2s60_burst_3_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_3_upstream_writedata = cpu_data_master_dbs_write_8;

  //byteaddress mux for std_2s60_burst_3/upstream, which is an e_mux
  assign std_2s60_burst_3_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_3_upstream = cpu_data_master_qualified_request_std_2s60_burst_3_upstream;

  //cpu/data_master saved-grant std_2s60_burst_3/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_3_upstream = cpu_data_master_requests_std_2s60_burst_3_upstream;

  //allow new arb cycle for std_2s60_burst_3/upstream, which is an e_assign
  assign std_2s60_burst_3_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_3_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_3_upstream_master_qreq_vector = 1;

  //std_2s60_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_3_upstream_firsttransfer = std_2s60_burst_3_upstream_begins_xfer ? std_2s60_burst_3_upstream_unreg_firsttransfer : std_2s60_burst_3_upstream_reg_firsttransfer;

  //std_2s60_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_3_upstream_unreg_firsttransfer = ~(std_2s60_burst_3_upstream_slavearbiterlockenable & std_2s60_burst_3_upstream_any_continuerequest);

  //std_2s60_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_3_upstream_begins_xfer)
          std_2s60_burst_3_upstream_reg_firsttransfer <= std_2s60_burst_3_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_3_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_3_upstream_next_bbt_burstcount = ((((std_2s60_burst_3_upstream_write) && (std_2s60_burst_3_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_3_upstream_burstcount - 1) :
    ((((std_2s60_burst_3_upstream_read) && (std_2s60_burst_3_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_3_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_3_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_3_upstream_begins_xfer)
          std_2s60_burst_3_upstream_bbt_burstcounter <= std_2s60_burst_3_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_3_upstream_beginbursttransfer_internal = std_2s60_burst_3_upstream_begins_xfer & (std_2s60_burst_3_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_3_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_3_upstream_read = cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_read;

  //std_2s60_burst_3_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_3_upstream_write = cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_write;

  //std_2s60_burst_3_upstream_address mux, which is an e_mux
  assign std_2s60_burst_3_upstream_address = {cpu_data_master_address_to_slave >> 2,
    cpu_data_master_dbs_address[1 : 0]};

  //d1_std_2s60_burst_3_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_3_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_3_upstream_end_xfer <= std_2s60_burst_3_upstream_end_xfer;
    end


  //std_2s60_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_3_upstream_waits_for_read = std_2s60_burst_3_upstream_in_a_read_cycle & std_2s60_burst_3_upstream_waitrequest_from_sa;

  //std_2s60_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_3_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_3_upstream_in_a_read_cycle;

  //std_2s60_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_3_upstream_waits_for_write = std_2s60_burst_3_upstream_in_a_write_cycle & std_2s60_burst_3_upstream_waitrequest_from_sa;

  //std_2s60_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_3_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_3_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_3_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_3_upstream_counter = 0;
  //std_2s60_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_3_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_3_upstream)? cpu_data_master_byteenable_std_2s60_burst_3_upstream :
    -1;

  assign {cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_3,
cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_2,
cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_1,
cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_0} = cpu_data_master_byteenable;
  assign cpu_data_master_byteenable_std_2s60_burst_3_upstream = ((cpu_data_master_dbs_address[1 : 0] == 0))? cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_0 :
    ((cpu_data_master_dbs_address[1 : 0] == 1))? cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_1 :
    ((cpu_data_master_dbs_address[1 : 0] == 2))? cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_2 :
    cpu_data_master_byteenable_std_2s60_burst_3_upstream_segment_3;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_3_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_3_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_3_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_3_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_3/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_3_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_3/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_3_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_flash_bus_avalon_slave_end_xfer,
                                                 ext_flash_s1_wait_counter_eq_0,
                                                 incoming_ext_flash_bus_data_with_Xs_converted_to_0,
                                                 reset_n,
                                                 std_2s60_burst_3_downstream_address,
                                                 std_2s60_burst_3_downstream_burstcount,
                                                 std_2s60_burst_3_downstream_byteenable,
                                                 std_2s60_burst_3_downstream_granted_ext_flash_s1,
                                                 std_2s60_burst_3_downstream_qualified_request_ext_flash_s1,
                                                 std_2s60_burst_3_downstream_read,
                                                 std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1,
                                                 std_2s60_burst_3_downstream_requests_ext_flash_s1,
                                                 std_2s60_burst_3_downstream_write,
                                                 std_2s60_burst_3_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_3_downstream_address_to_slave,
                                                 std_2s60_burst_3_downstream_latency_counter,
                                                 std_2s60_burst_3_downstream_readdata,
                                                 std_2s60_burst_3_downstream_readdatavalid,
                                                 std_2s60_burst_3_downstream_reset_n,
                                                 std_2s60_burst_3_downstream_waitrequest
                                              )
;

  output  [ 23: 0] std_2s60_burst_3_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_3_downstream_latency_counter;
  output  [  7: 0] std_2s60_burst_3_downstream_readdata;
  output           std_2s60_burst_3_downstream_readdatavalid;
  output           std_2s60_burst_3_downstream_reset_n;
  output           std_2s60_burst_3_downstream_waitrequest;
  input            clk;
  input            d1_ext_flash_bus_avalon_slave_end_xfer;
  input            ext_flash_s1_wait_counter_eq_0;
  input   [  7: 0] incoming_ext_flash_bus_data_with_Xs_converted_to_0;
  input            reset_n;
  input   [ 23: 0] std_2s60_burst_3_downstream_address;
  input            std_2s60_burst_3_downstream_burstcount;
  input            std_2s60_burst_3_downstream_byteenable;
  input            std_2s60_burst_3_downstream_granted_ext_flash_s1;
  input            std_2s60_burst_3_downstream_qualified_request_ext_flash_s1;
  input            std_2s60_burst_3_downstream_read;
  input            std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1;
  input            std_2s60_burst_3_downstream_requests_ext_flash_s1;
  input            std_2s60_burst_3_downstream_write;
  input   [  7: 0] std_2s60_burst_3_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_3_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_3_downstream_readdatavalid;
  wire             r_0;
  reg     [ 23: 0] std_2s60_burst_3_downstream_address_last_time;
  wire    [ 23: 0] std_2s60_burst_3_downstream_address_to_slave;
  reg              std_2s60_burst_3_downstream_burstcount_last_time;
  reg              std_2s60_burst_3_downstream_byteenable_last_time;
  wire             std_2s60_burst_3_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_3_downstream_latency_counter;
  reg              std_2s60_burst_3_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_3_downstream_read_last_time;
  wire    [  7: 0] std_2s60_burst_3_downstream_readdata;
  wire             std_2s60_burst_3_downstream_readdatavalid;
  wire             std_2s60_burst_3_downstream_reset_n;
  wire             std_2s60_burst_3_downstream_run;
  wire             std_2s60_burst_3_downstream_waitrequest;
  reg              std_2s60_burst_3_downstream_write_last_time;
  reg     [  7: 0] std_2s60_burst_3_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_3_downstream_requests_ext_flash_s1) & (std_2s60_burst_3_downstream_granted_ext_flash_s1 | ~std_2s60_burst_3_downstream_qualified_request_ext_flash_s1) & ((~std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_3_downstream_read | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_ext_flash_bus_avalon_slave_end_xfer)) & std_2s60_burst_3_downstream_read))) & ((~std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 | ~std_2s60_burst_3_downstream_write | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_ext_flash_bus_avalon_slave_end_xfer)) & std_2s60_burst_3_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_3_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_3_downstream_address_to_slave = std_2s60_burst_3_downstream_address;

  //std_2s60_burst_3_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_3_downstream_read_but_no_slave_selected <= std_2s60_burst_3_downstream_read & std_2s60_burst_3_downstream_run & ~std_2s60_burst_3_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_3_downstream_is_granted_some_slave = std_2s60_burst_3_downstream_granted_ext_flash_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_3_downstream_readdatavalid = std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_3_downstream_readdatavalid = std_2s60_burst_3_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_3_downstream_readdatavalid;

  //std_2s60_burst_3/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_3_downstream_readdata = incoming_ext_flash_bus_data_with_Xs_converted_to_0;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_3_downstream_waitrequest = ~std_2s60_burst_3_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_3_downstream_latency_counter <= p1_std_2s60_burst_3_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_3_downstream_latency_counter = ((std_2s60_burst_3_downstream_run & std_2s60_burst_3_downstream_read))? latency_load_value :
    (std_2s60_burst_3_downstream_latency_counter)? std_2s60_burst_3_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {2 {std_2s60_burst_3_downstream_requests_ext_flash_s1}} & 2;

  //std_2s60_burst_3_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_3_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_3_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_address_last_time <= std_2s60_burst_3_downstream_address;
    end


  //std_2s60_burst_3/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_3_downstream_waitrequest & (std_2s60_burst_3_downstream_read | std_2s60_burst_3_downstream_write);
    end


  //std_2s60_burst_3_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_address != std_2s60_burst_3_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_3_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_burstcount_last_time <= std_2s60_burst_3_downstream_burstcount;
    end


  //std_2s60_burst_3_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_burstcount != std_2s60_burst_3_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_3_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_byteenable_last_time <= std_2s60_burst_3_downstream_byteenable;
    end


  //std_2s60_burst_3_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_byteenable != std_2s60_burst_3_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_3_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_read_last_time <= std_2s60_burst_3_downstream_read;
    end


  //std_2s60_burst_3_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_read != std_2s60_burst_3_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_3_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_write_last_time <= std_2s60_burst_3_downstream_write;
    end


  //std_2s60_burst_3_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_write != std_2s60_burst_3_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_3_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_3_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_3_downstream_writedata_last_time <= std_2s60_burst_3_downstream_writedata;
    end


  //std_2s60_burst_3_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_3_downstream_writedata != std_2s60_burst_3_downstream_writedata_last_time) & std_2s60_burst_3_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_3_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_4_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_4_upstream_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_4_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_instruction_master_address_to_slave,
                                               cpu_instruction_master_burstcount,
                                               cpu_instruction_master_latency_counter,
                                               cpu_instruction_master_read,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                               reset_n,
                                               std_2s60_burst_4_upstream_readdata,
                                               std_2s60_burst_4_upstream_readdatavalid,
                                               std_2s60_burst_4_upstream_waitrequest,

                                              // outputs:
                                               cpu_instruction_master_granted_std_2s60_burst_4_upstream,
                                               cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                               cpu_instruction_master_requests_std_2s60_burst_4_upstream,
                                               d1_std_2s60_burst_4_upstream_end_xfer,
                                               std_2s60_burst_4_upstream_address,
                                               std_2s60_burst_4_upstream_byteaddress,
                                               std_2s60_burst_4_upstream_byteenable,
                                               std_2s60_burst_4_upstream_debugaccess,
                                               std_2s60_burst_4_upstream_read,
                                               std_2s60_burst_4_upstream_readdata_from_sa,
                                               std_2s60_burst_4_upstream_waitrequest_from_sa,
                                               std_2s60_burst_4_upstream_write
                                            )
;

  output           cpu_instruction_master_granted_std_2s60_burst_4_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_4_upstream;
  output           d1_std_2s60_burst_4_upstream_end_xfer;
  output  [ 19: 0] std_2s60_burst_4_upstream_address;
  output  [ 21: 0] std_2s60_burst_4_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_4_upstream_byteenable;
  output           std_2s60_burst_4_upstream_debugaccess;
  output           std_2s60_burst_4_upstream_read;
  output  [ 31: 0] std_2s60_burst_4_upstream_readdata_from_sa;
  output           std_2s60_burst_4_upstream_waitrequest_from_sa;
  output           std_2s60_burst_4_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_4_upstream_readdata;
  input            std_2s60_burst_4_upstream_readdatavalid;
  input            std_2s60_burst_4_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_4_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_4_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_4_upstream_load_fifo;
  wire    [ 19: 0] std_2s60_burst_4_upstream_address;
  wire             std_2s60_burst_4_upstream_allgrants;
  wire             std_2s60_burst_4_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_4_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_4_upstream_any_continuerequest;
  wire             std_2s60_burst_4_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_4_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_4_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_4_upstream_arb_share_set_values;
  wire             std_2s60_burst_4_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_4_upstream_begins_xfer;
  wire             std_2s60_burst_4_upstream_burstcount_fifo_empty;
  wire    [ 21: 0] std_2s60_burst_4_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_4_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_4_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_4_upstream_current_burst_minus_one;
  wire             std_2s60_burst_4_upstream_debugaccess;
  wire             std_2s60_burst_4_upstream_end_xfer;
  wire             std_2s60_burst_4_upstream_firsttransfer;
  wire             std_2s60_burst_4_upstream_grant_vector;
  wire             std_2s60_burst_4_upstream_in_a_read_cycle;
  wire             std_2s60_burst_4_upstream_in_a_write_cycle;
  reg              std_2s60_burst_4_upstream_load_fifo;
  wire             std_2s60_burst_4_upstream_master_qreq_vector;
  wire             std_2s60_burst_4_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_4_upstream_next_burst_count;
  wire             std_2s60_burst_4_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_4_upstream_read;
  wire    [ 31: 0] std_2s60_burst_4_upstream_readdata_from_sa;
  wire             std_2s60_burst_4_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_4_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_4_upstream_selected_burstcount;
  reg              std_2s60_burst_4_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_4_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_4_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_4_upstream_transaction_burst_count;
  wire             std_2s60_burst_4_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_4_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_4_upstream_waits_for_read;
  wire             std_2s60_burst_4_upstream_waits_for_write;
  wire             std_2s60_burst_4_upstream_write;
  wire             wait_for_std_2s60_burst_4_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_4_upstream_end_xfer;
    end


  assign std_2s60_burst_4_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream));
  //assign std_2s60_burst_4_upstream_readdatavalid_from_sa = std_2s60_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_4_upstream_readdatavalid_from_sa = std_2s60_burst_4_upstream_readdatavalid;

  //assign std_2s60_burst_4_upstream_readdata_from_sa = std_2s60_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_4_upstream_readdata_from_sa = std_2s60_burst_4_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_4_upstream = (({cpu_instruction_master_address_to_slave[25 : 20] , 20'b0} == 26'h2200000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_4_upstream_waitrequest_from_sa = std_2s60_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_4_upstream_waitrequest_from_sa = std_2s60_burst_4_upstream_waitrequest;

  //std_2s60_burst_4_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_4_upstream_arb_share_set_values = 1;

  //std_2s60_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_4_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_4_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_4_upstream;

  //std_2s60_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_4_upstream_arb_share_counter_next_value = std_2s60_burst_4_upstream_firsttransfer ? (std_2s60_burst_4_upstream_arb_share_set_values - 1) : |std_2s60_burst_4_upstream_arb_share_counter ? (std_2s60_burst_4_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_4_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_4_upstream_allgrants = |std_2s60_burst_4_upstream_grant_vector;

  //std_2s60_burst_4_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_4_upstream_end_xfer = ~(std_2s60_burst_4_upstream_waits_for_read | std_2s60_burst_4_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream = std_2s60_burst_4_upstream_end_xfer & (~std_2s60_burst_4_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_4_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream & std_2s60_burst_4_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream & ~std_2s60_burst_4_upstream_non_bursting_master_requests);

  //std_2s60_burst_4_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_4_upstream_arb_counter_enable)
          std_2s60_burst_4_upstream_arb_share_counter <= std_2s60_burst_4_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_4_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_4_upstream & ~std_2s60_burst_4_upstream_non_bursting_master_requests))
          std_2s60_burst_4_upstream_slavearbiterlockenable <= |std_2s60_burst_4_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_4/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_4_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_4_upstream_slavearbiterlockenable2 = |std_2s60_burst_4_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_4/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_4_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_4_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream = cpu_instruction_master_requests_std_2s60_burst_4_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_4_upstream_move_on_to_next_transaction = std_2s60_burst_4_upstream_this_cycle_is_the_last_burst & std_2s60_burst_4_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_4_upstream, which is an e_mux
  assign std_2s60_burst_4_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_4_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_4_upstream_module burstcount_fifo_for_std_2s60_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_4_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_4_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_4_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_4_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read & std_2s60_burst_4_upstream_load_fifo & ~(std_2s60_burst_4_upstream_this_cycle_is_the_last_burst & std_2s60_burst_4_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_4_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_4_upstream_current_burst_minus_one = std_2s60_burst_4_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_4_upstream, which is an e_mux
  assign std_2s60_burst_4_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read) & ~std_2s60_burst_4_upstream_load_fifo))? std_2s60_burst_4_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read & std_2s60_burst_4_upstream_this_cycle_is_the_last_burst & std_2s60_burst_4_upstream_burstcount_fifo_empty))? std_2s60_burst_4_upstream_selected_burstcount :
    (std_2s60_burst_4_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_4_upstream_transaction_burst_count :
    std_2s60_burst_4_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_4_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_upstream_current_burst <= 0;
      else if (std_2s60_burst_4_upstream_readdatavalid_from_sa | (~std_2s60_burst_4_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read)))
          std_2s60_burst_4_upstream_current_burst <= std_2s60_burst_4_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_4_upstream_load_fifo = (~std_2s60_burst_4_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read) & std_2s60_burst_4_upstream_load_fifo))? 1 :
    ~std_2s60_burst_4_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read) & ~std_2s60_burst_4_upstream_load_fifo | std_2s60_burst_4_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_4_upstream_load_fifo <= p0_std_2s60_burst_4_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_4_upstream, which is an e_assign
  assign std_2s60_burst_4_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_4_upstream_current_burst_minus_one) & std_2s60_burst_4_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_4_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_4_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_4_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_4_upstream),
      .full                 (),
      .read                 (std_2s60_burst_4_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_4_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_4_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream = std_2s60_burst_4_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_4/upstream, which is an e_mux
  assign std_2s60_burst_4_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_4_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_4/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_4_upstream = cpu_instruction_master_requests_std_2s60_burst_4_upstream;

  //allow new arb cycle for std_2s60_burst_4/upstream, which is an e_assign
  assign std_2s60_burst_4_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_4_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_4_upstream_master_qreq_vector = 1;

  //std_2s60_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_4_upstream_firsttransfer = std_2s60_burst_4_upstream_begins_xfer ? std_2s60_burst_4_upstream_unreg_firsttransfer : std_2s60_burst_4_upstream_reg_firsttransfer;

  //std_2s60_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_4_upstream_unreg_firsttransfer = ~(std_2s60_burst_4_upstream_slavearbiterlockenable & std_2s60_burst_4_upstream_any_continuerequest);

  //std_2s60_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_4_upstream_begins_xfer)
          std_2s60_burst_4_upstream_reg_firsttransfer <= std_2s60_burst_4_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_4_upstream_beginbursttransfer_internal = std_2s60_burst_4_upstream_begins_xfer;

  //std_2s60_burst_4_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_4_upstream_read = cpu_instruction_master_granted_std_2s60_burst_4_upstream & cpu_instruction_master_read;

  //std_2s60_burst_4_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_4_upstream_write = 0;

  //std_2s60_burst_4_upstream_address mux, which is an e_mux
  assign std_2s60_burst_4_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_std_2s60_burst_4_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_4_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_4_upstream_end_xfer <= std_2s60_burst_4_upstream_end_xfer;
    end


  //std_2s60_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_4_upstream_waits_for_read = std_2s60_burst_4_upstream_in_a_read_cycle & std_2s60_burst_4_upstream_waitrequest_from_sa;

  //std_2s60_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_4_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_4_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_4_upstream_in_a_read_cycle;

  //std_2s60_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_4_upstream_waits_for_write = std_2s60_burst_4_upstream_in_a_write_cycle & std_2s60_burst_4_upstream_waitrequest_from_sa;

  //std_2s60_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_4_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_4_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_4_upstream_counter = 0;
  //std_2s60_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_4_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_4_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_4/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_4_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_4/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_4_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_ram_bus_avalon_slave_end_xfer,
                                                 ext_ram_s1_wait_counter_eq_0,
                                                 incoming_ext_ram_bus_data,
                                                 lan91c111_s1_wait_counter_eq_0,
                                                 reset_n,
                                                 std_2s60_burst_4_downstream_address,
                                                 std_2s60_burst_4_downstream_burstcount,
                                                 std_2s60_burst_4_downstream_byteenable,
                                                 std_2s60_burst_4_downstream_granted_ext_ram_s1,
                                                 std_2s60_burst_4_downstream_granted_lan91c111_s1,
                                                 std_2s60_burst_4_downstream_qualified_request_ext_ram_s1,
                                                 std_2s60_burst_4_downstream_qualified_request_lan91c111_s1,
                                                 std_2s60_burst_4_downstream_read,
                                                 std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1,
                                                 std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1,
                                                 std_2s60_burst_4_downstream_requests_ext_ram_s1,
                                                 std_2s60_burst_4_downstream_requests_lan91c111_s1,
                                                 std_2s60_burst_4_downstream_write,
                                                 std_2s60_burst_4_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_4_downstream_address_to_slave,
                                                 std_2s60_burst_4_downstream_latency_counter,
                                                 std_2s60_burst_4_downstream_readdata,
                                                 std_2s60_burst_4_downstream_readdatavalid,
                                                 std_2s60_burst_4_downstream_reset_n,
                                                 std_2s60_burst_4_downstream_waitrequest
                                              )
;

  output  [ 19: 0] std_2s60_burst_4_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_4_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_4_downstream_readdata;
  output           std_2s60_burst_4_downstream_readdatavalid;
  output           std_2s60_burst_4_downstream_reset_n;
  output           std_2s60_burst_4_downstream_waitrequest;
  input            clk;
  input            d1_ext_ram_bus_avalon_slave_end_xfer;
  input            ext_ram_s1_wait_counter_eq_0;
  input   [ 31: 0] incoming_ext_ram_bus_data;
  input            lan91c111_s1_wait_counter_eq_0;
  input            reset_n;
  input   [ 19: 0] std_2s60_burst_4_downstream_address;
  input            std_2s60_burst_4_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_4_downstream_byteenable;
  input            std_2s60_burst_4_downstream_granted_ext_ram_s1;
  input            std_2s60_burst_4_downstream_granted_lan91c111_s1;
  input            std_2s60_burst_4_downstream_qualified_request_ext_ram_s1;
  input            std_2s60_burst_4_downstream_qualified_request_lan91c111_s1;
  input            std_2s60_burst_4_downstream_read;
  input            std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1;
  input            std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1;
  input            std_2s60_burst_4_downstream_requests_ext_ram_s1;
  input            std_2s60_burst_4_downstream_requests_lan91c111_s1;
  input            std_2s60_burst_4_downstream_write;
  input   [ 31: 0] std_2s60_burst_4_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_4_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_4_downstream_readdatavalid;
  wire             r_0;
  reg     [ 19: 0] std_2s60_burst_4_downstream_address_last_time;
  wire    [ 19: 0] std_2s60_burst_4_downstream_address_to_slave;
  reg              std_2s60_burst_4_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_4_downstream_byteenable_last_time;
  wire             std_2s60_burst_4_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_4_downstream_latency_counter;
  reg              std_2s60_burst_4_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_4_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_4_downstream_readdata;
  wire             std_2s60_burst_4_downstream_readdatavalid;
  wire             std_2s60_burst_4_downstream_reset_n;
  wire             std_2s60_burst_4_downstream_run;
  wire             std_2s60_burst_4_downstream_waitrequest;
  reg              std_2s60_burst_4_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_4_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_4_downstream_requests_lan91c111_s1) & (std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_4_downstream_requests_ext_ram_s1) & (std_2s60_burst_4_downstream_granted_lan91c111_s1 | ~std_2s60_burst_4_downstream_qualified_request_lan91c111_s1) & (std_2s60_burst_4_downstream_granted_ext_ram_s1 | ~std_2s60_burst_4_downstream_qualified_request_ext_ram_s1) & ((~std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_4_downstream_read | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_4_downstream_read))) & ((~std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_4_downstream_write | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_4_downstream_write))) & ((~std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_4_downstream_read | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_4_downstream_read))) & ((~std_2s60_burst_4_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_4_downstream_write | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_4_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_4_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_4_downstream_address_to_slave = std_2s60_burst_4_downstream_address;

  //std_2s60_burst_4_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_4_downstream_read_but_no_slave_selected <= std_2s60_burst_4_downstream_read & std_2s60_burst_4_downstream_run & ~std_2s60_burst_4_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_4_downstream_is_granted_some_slave = std_2s60_burst_4_downstream_granted_lan91c111_s1 |
    std_2s60_burst_4_downstream_granted_ext_ram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_4_downstream_readdatavalid = std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1 |
    std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_4_downstream_readdatavalid = std_2s60_burst_4_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_4_downstream_readdatavalid |
    std_2s60_burst_4_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_4_downstream_readdatavalid;

  //std_2s60_burst_4/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_4_downstream_readdata = ({32 {~std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1}} | incoming_ext_ram_bus_data) &
    ({32 {~std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1}} | incoming_ext_ram_bus_data);

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_4_downstream_waitrequest = ~std_2s60_burst_4_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_4_downstream_latency_counter <= p1_std_2s60_burst_4_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_4_downstream_latency_counter = ((std_2s60_burst_4_downstream_run & std_2s60_burst_4_downstream_read))? latency_load_value :
    (std_2s60_burst_4_downstream_latency_counter)? std_2s60_burst_4_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {std_2s60_burst_4_downstream_requests_lan91c111_s1}} & 2) |
    ({2 {std_2s60_burst_4_downstream_requests_ext_ram_s1}} & 2);

  //std_2s60_burst_4_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_4_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_4_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_address_last_time <= std_2s60_burst_4_downstream_address;
    end


  //std_2s60_burst_4/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_4_downstream_waitrequest & (std_2s60_burst_4_downstream_read | std_2s60_burst_4_downstream_write);
    end


  //std_2s60_burst_4_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_address != std_2s60_burst_4_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_4_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_burstcount_last_time <= std_2s60_burst_4_downstream_burstcount;
    end


  //std_2s60_burst_4_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_burstcount != std_2s60_burst_4_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_4_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_byteenable_last_time <= std_2s60_burst_4_downstream_byteenable;
    end


  //std_2s60_burst_4_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_byteenable != std_2s60_burst_4_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_4_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_read_last_time <= std_2s60_burst_4_downstream_read;
    end


  //std_2s60_burst_4_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_read != std_2s60_burst_4_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_4_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_write_last_time <= std_2s60_burst_4_downstream_write;
    end


  //std_2s60_burst_4_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_write != std_2s60_burst_4_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_4_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_4_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_4_downstream_writedata_last_time <= std_2s60_burst_4_downstream_writedata;
    end


  //std_2s60_burst_4_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_4_downstream_writedata != std_2s60_burst_4_downstream_writedata_last_time) & std_2s60_burst_4_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_4_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_5_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_5_upstream_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_5_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_burstcount,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_debugaccess,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                               cpu_data_master_write,
                                               cpu_data_master_writedata,
                                               reset_n,
                                               std_2s60_burst_5_upstream_readdata,
                                               std_2s60_burst_5_upstream_readdatavalid,
                                               std_2s60_burst_5_upstream_waitrequest,

                                              // outputs:
                                               cpu_data_master_granted_std_2s60_burst_5_upstream,
                                               cpu_data_master_qualified_request_std_2s60_burst_5_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                               cpu_data_master_requests_std_2s60_burst_5_upstream,
                                               d1_std_2s60_burst_5_upstream_end_xfer,
                                               std_2s60_burst_5_upstream_address,
                                               std_2s60_burst_5_upstream_burstcount,
                                               std_2s60_burst_5_upstream_byteaddress,
                                               std_2s60_burst_5_upstream_byteenable,
                                               std_2s60_burst_5_upstream_debugaccess,
                                               std_2s60_burst_5_upstream_read,
                                               std_2s60_burst_5_upstream_readdata_from_sa,
                                               std_2s60_burst_5_upstream_waitrequest_from_sa,
                                               std_2s60_burst_5_upstream_write,
                                               std_2s60_burst_5_upstream_writedata
                                            )
;

  output           cpu_data_master_granted_std_2s60_burst_5_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_5_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_5_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_5_upstream;
  output           d1_std_2s60_burst_5_upstream_end_xfer;
  output  [ 19: 0] std_2s60_burst_5_upstream_address;
  output  [  3: 0] std_2s60_burst_5_upstream_burstcount;
  output  [ 21: 0] std_2s60_burst_5_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_5_upstream_byteenable;
  output           std_2s60_burst_5_upstream_debugaccess;
  output           std_2s60_burst_5_upstream_read;
  output  [ 31: 0] std_2s60_burst_5_upstream_readdata_from_sa;
  output           std_2s60_burst_5_upstream_waitrequest_from_sa;
  output           std_2s60_burst_5_upstream_write;
  output  [ 31: 0] std_2s60_burst_5_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_5_upstream_readdata;
  input            std_2s60_burst_5_upstream_readdatavalid;
  input            std_2s60_burst_5_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_5_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_5_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_5_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_5_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_5_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_5_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_5_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_5_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_5_upstream_load_fifo;
  wire    [ 19: 0] std_2s60_burst_5_upstream_address;
  wire             std_2s60_burst_5_upstream_allgrants;
  wire             std_2s60_burst_5_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_5_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_5_upstream_any_continuerequest;
  wire             std_2s60_burst_5_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_5_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_5_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_5_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_5_upstream_bbt_burstcounter;
  wire             std_2s60_burst_5_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_5_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_5_upstream_burstcount;
  wire             std_2s60_burst_5_upstream_burstcount_fifo_empty;
  wire    [ 21: 0] std_2s60_burst_5_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_5_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_5_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_5_upstream_current_burst_minus_one;
  wire             std_2s60_burst_5_upstream_debugaccess;
  wire             std_2s60_burst_5_upstream_end_xfer;
  wire             std_2s60_burst_5_upstream_firsttransfer;
  wire             std_2s60_burst_5_upstream_grant_vector;
  wire             std_2s60_burst_5_upstream_in_a_read_cycle;
  wire             std_2s60_burst_5_upstream_in_a_write_cycle;
  reg              std_2s60_burst_5_upstream_load_fifo;
  wire             std_2s60_burst_5_upstream_master_qreq_vector;
  wire             std_2s60_burst_5_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_5_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_5_upstream_next_burst_count;
  wire             std_2s60_burst_5_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_5_upstream_read;
  wire    [ 31: 0] std_2s60_burst_5_upstream_readdata_from_sa;
  wire             std_2s60_burst_5_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_5_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_5_upstream_selected_burstcount;
  reg              std_2s60_burst_5_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_5_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_5_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_5_upstream_transaction_burst_count;
  wire             std_2s60_burst_5_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_5_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_5_upstream_waits_for_read;
  wire             std_2s60_burst_5_upstream_waits_for_write;
  wire             std_2s60_burst_5_upstream_write;
  wire    [ 31: 0] std_2s60_burst_5_upstream_writedata;
  wire             wait_for_std_2s60_burst_5_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_5_upstream_end_xfer;
    end


  assign std_2s60_burst_5_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_5_upstream));
  //assign std_2s60_burst_5_upstream_readdatavalid_from_sa = std_2s60_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_5_upstream_readdatavalid_from_sa = std_2s60_burst_5_upstream_readdatavalid;

  //assign std_2s60_burst_5_upstream_readdata_from_sa = std_2s60_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_5_upstream_readdata_from_sa = std_2s60_burst_5_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_5_upstream = ({cpu_data_master_address_to_slave[25 : 20] , 20'b0} == 26'h2200000) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_5_upstream_waitrequest_from_sa = std_2s60_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_5_upstream_waitrequest_from_sa = std_2s60_burst_5_upstream_waitrequest;

  //std_2s60_burst_5_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_5_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_5_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_5_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_5_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_5_upstream;

  //std_2s60_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_5_upstream_arb_share_counter_next_value = std_2s60_burst_5_upstream_firsttransfer ? (std_2s60_burst_5_upstream_arb_share_set_values - 1) : |std_2s60_burst_5_upstream_arb_share_counter ? (std_2s60_burst_5_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_5_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_5_upstream_allgrants = |std_2s60_burst_5_upstream_grant_vector;

  //std_2s60_burst_5_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_5_upstream_end_xfer = ~(std_2s60_burst_5_upstream_waits_for_read | std_2s60_burst_5_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream = std_2s60_burst_5_upstream_end_xfer & (~std_2s60_burst_5_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_5_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream & std_2s60_burst_5_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream & ~std_2s60_burst_5_upstream_non_bursting_master_requests);

  //std_2s60_burst_5_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_5_upstream_arb_counter_enable)
          std_2s60_burst_5_upstream_arb_share_counter <= std_2s60_burst_5_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_5_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_5_upstream & ~std_2s60_burst_5_upstream_non_bursting_master_requests))
          std_2s60_burst_5_upstream_slavearbiterlockenable <= |std_2s60_burst_5_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_5/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_5_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_5_upstream_slavearbiterlockenable2 = |std_2s60_burst_5_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_5/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_5_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_5_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_5_upstream = cpu_data_master_requests_std_2s60_burst_5_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_5_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_5_upstream_move_on_to_next_transaction = std_2s60_burst_5_upstream_this_cycle_is_the_last_burst & std_2s60_burst_5_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_5_upstream, which is an e_mux
  assign std_2s60_burst_5_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_5_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_5_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_5_upstream_module burstcount_fifo_for_std_2s60_burst_5_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_5_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_5_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_5_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_5_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read & std_2s60_burst_5_upstream_load_fifo & ~(std_2s60_burst_5_upstream_this_cycle_is_the_last_burst & std_2s60_burst_5_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_5_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_5_upstream_current_burst_minus_one = std_2s60_burst_5_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_5_upstream, which is an e_mux
  assign std_2s60_burst_5_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read) & ~std_2s60_burst_5_upstream_load_fifo))? std_2s60_burst_5_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read & std_2s60_burst_5_upstream_this_cycle_is_the_last_burst & std_2s60_burst_5_upstream_burstcount_fifo_empty))? std_2s60_burst_5_upstream_selected_burstcount :
    (std_2s60_burst_5_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_5_upstream_transaction_burst_count :
    std_2s60_burst_5_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_5_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_current_burst <= 0;
      else if (std_2s60_burst_5_upstream_readdatavalid_from_sa | (~std_2s60_burst_5_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read)))
          std_2s60_burst_5_upstream_current_burst <= std_2s60_burst_5_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_5_upstream_load_fifo = (~std_2s60_burst_5_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read) & std_2s60_burst_5_upstream_load_fifo))? 1 :
    ~std_2s60_burst_5_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read) & ~std_2s60_burst_5_upstream_load_fifo | std_2s60_burst_5_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_5_upstream_load_fifo <= p0_std_2s60_burst_5_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_5_upstream, which is an e_assign
  assign std_2s60_burst_5_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_5_upstream_current_burst_minus_one) & std_2s60_burst_5_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_5_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_5_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_5_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_5_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_5_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_5_upstream),
      .full                 (),
      .read                 (std_2s60_burst_5_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_5_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_5_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_5_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_5_upstream = std_2s60_burst_5_upstream_readdatavalid_from_sa;

  //std_2s60_burst_5_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_5_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_5/upstream, which is an e_mux
  assign std_2s60_burst_5_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_5_upstream = cpu_data_master_qualified_request_std_2s60_burst_5_upstream;

  //cpu/data_master saved-grant std_2s60_burst_5/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_5_upstream = cpu_data_master_requests_std_2s60_burst_5_upstream;

  //allow new arb cycle for std_2s60_burst_5/upstream, which is an e_assign
  assign std_2s60_burst_5_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_5_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_5_upstream_master_qreq_vector = 1;

  //std_2s60_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_5_upstream_firsttransfer = std_2s60_burst_5_upstream_begins_xfer ? std_2s60_burst_5_upstream_unreg_firsttransfer : std_2s60_burst_5_upstream_reg_firsttransfer;

  //std_2s60_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_5_upstream_unreg_firsttransfer = ~(std_2s60_burst_5_upstream_slavearbiterlockenable & std_2s60_burst_5_upstream_any_continuerequest);

  //std_2s60_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_5_upstream_begins_xfer)
          std_2s60_burst_5_upstream_reg_firsttransfer <= std_2s60_burst_5_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_5_upstream_next_bbt_burstcount = ((((std_2s60_burst_5_upstream_write) && (std_2s60_burst_5_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_5_upstream_burstcount - 1) :
    ((((std_2s60_burst_5_upstream_read) && (std_2s60_burst_5_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_5_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_5_upstream_begins_xfer)
          std_2s60_burst_5_upstream_bbt_burstcounter <= std_2s60_burst_5_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_5_upstream_beginbursttransfer_internal = std_2s60_burst_5_upstream_begins_xfer & (std_2s60_burst_5_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_5_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_5_upstream_read = cpu_data_master_granted_std_2s60_burst_5_upstream & cpu_data_master_read;

  //std_2s60_burst_5_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_5_upstream_write = cpu_data_master_granted_std_2s60_burst_5_upstream & cpu_data_master_write;

  //std_2s60_burst_5_upstream_address mux, which is an e_mux
  assign std_2s60_burst_5_upstream_address = cpu_data_master_address_to_slave;

  //d1_std_2s60_burst_5_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_5_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_5_upstream_end_xfer <= std_2s60_burst_5_upstream_end_xfer;
    end


  //std_2s60_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_5_upstream_waits_for_read = std_2s60_burst_5_upstream_in_a_read_cycle & std_2s60_burst_5_upstream_waitrequest_from_sa;

  //std_2s60_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_5_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_5_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_5_upstream_in_a_read_cycle;

  //std_2s60_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_5_upstream_waits_for_write = std_2s60_burst_5_upstream_in_a_write_cycle & std_2s60_burst_5_upstream_waitrequest_from_sa;

  //std_2s60_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_5_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_5_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_5_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_5_upstream_counter = 0;
  //std_2s60_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_5_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_5_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_5_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_5_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_5_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_5_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_5/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_5_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_5/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_5_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_ram_bus_avalon_slave_end_xfer,
                                                 ext_ram_s1_wait_counter_eq_0,
                                                 incoming_ext_ram_bus_data,
                                                 lan91c111_s1_wait_counter_eq_0,
                                                 reset_n,
                                                 std_2s60_burst_5_downstream_address,
                                                 std_2s60_burst_5_downstream_burstcount,
                                                 std_2s60_burst_5_downstream_byteenable,
                                                 std_2s60_burst_5_downstream_granted_ext_ram_s1,
                                                 std_2s60_burst_5_downstream_granted_lan91c111_s1,
                                                 std_2s60_burst_5_downstream_qualified_request_ext_ram_s1,
                                                 std_2s60_burst_5_downstream_qualified_request_lan91c111_s1,
                                                 std_2s60_burst_5_downstream_read,
                                                 std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1,
                                                 std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1,
                                                 std_2s60_burst_5_downstream_requests_ext_ram_s1,
                                                 std_2s60_burst_5_downstream_requests_lan91c111_s1,
                                                 std_2s60_burst_5_downstream_write,
                                                 std_2s60_burst_5_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_5_downstream_address_to_slave,
                                                 std_2s60_burst_5_downstream_latency_counter,
                                                 std_2s60_burst_5_downstream_readdata,
                                                 std_2s60_burst_5_downstream_readdatavalid,
                                                 std_2s60_burst_5_downstream_reset_n,
                                                 std_2s60_burst_5_downstream_waitrequest
                                              )
;

  output  [ 19: 0] std_2s60_burst_5_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_5_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_5_downstream_readdata;
  output           std_2s60_burst_5_downstream_readdatavalid;
  output           std_2s60_burst_5_downstream_reset_n;
  output           std_2s60_burst_5_downstream_waitrequest;
  input            clk;
  input            d1_ext_ram_bus_avalon_slave_end_xfer;
  input            ext_ram_s1_wait_counter_eq_0;
  input   [ 31: 0] incoming_ext_ram_bus_data;
  input            lan91c111_s1_wait_counter_eq_0;
  input            reset_n;
  input   [ 19: 0] std_2s60_burst_5_downstream_address;
  input            std_2s60_burst_5_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_5_downstream_byteenable;
  input            std_2s60_burst_5_downstream_granted_ext_ram_s1;
  input            std_2s60_burst_5_downstream_granted_lan91c111_s1;
  input            std_2s60_burst_5_downstream_qualified_request_ext_ram_s1;
  input            std_2s60_burst_5_downstream_qualified_request_lan91c111_s1;
  input            std_2s60_burst_5_downstream_read;
  input            std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1;
  input            std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1;
  input            std_2s60_burst_5_downstream_requests_ext_ram_s1;
  input            std_2s60_burst_5_downstream_requests_lan91c111_s1;
  input            std_2s60_burst_5_downstream_write;
  input   [ 31: 0] std_2s60_burst_5_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_5_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_5_downstream_readdatavalid;
  wire             r_0;
  reg     [ 19: 0] std_2s60_burst_5_downstream_address_last_time;
  wire    [ 19: 0] std_2s60_burst_5_downstream_address_to_slave;
  reg              std_2s60_burst_5_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_5_downstream_byteenable_last_time;
  wire             std_2s60_burst_5_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_5_downstream_latency_counter;
  reg              std_2s60_burst_5_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_5_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_5_downstream_readdata;
  wire             std_2s60_burst_5_downstream_readdatavalid;
  wire             std_2s60_burst_5_downstream_reset_n;
  wire             std_2s60_burst_5_downstream_run;
  wire             std_2s60_burst_5_downstream_waitrequest;
  reg              std_2s60_burst_5_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_5_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_5_downstream_requests_lan91c111_s1) & (std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_5_downstream_requests_ext_ram_s1) & (std_2s60_burst_5_downstream_granted_lan91c111_s1 | ~std_2s60_burst_5_downstream_qualified_request_lan91c111_s1) & (std_2s60_burst_5_downstream_granted_ext_ram_s1 | ~std_2s60_burst_5_downstream_qualified_request_ext_ram_s1) & ((~std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_5_downstream_read | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_5_downstream_read))) & ((~std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_5_downstream_write | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_5_downstream_write))) & ((~std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_5_downstream_read | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_5_downstream_read))) & ((~std_2s60_burst_5_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_5_downstream_write | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_5_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_5_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_5_downstream_address_to_slave = std_2s60_burst_5_downstream_address;

  //std_2s60_burst_5_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_5_downstream_read_but_no_slave_selected <= std_2s60_burst_5_downstream_read & std_2s60_burst_5_downstream_run & ~std_2s60_burst_5_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_5_downstream_is_granted_some_slave = std_2s60_burst_5_downstream_granted_lan91c111_s1 |
    std_2s60_burst_5_downstream_granted_ext_ram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_5_downstream_readdatavalid = std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1 |
    std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_5_downstream_readdatavalid = std_2s60_burst_5_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_5_downstream_readdatavalid |
    std_2s60_burst_5_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_5_downstream_readdatavalid;

  //std_2s60_burst_5/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_5_downstream_readdata = ({32 {~std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1}} | incoming_ext_ram_bus_data) &
    ({32 {~std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1}} | incoming_ext_ram_bus_data);

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_5_downstream_waitrequest = ~std_2s60_burst_5_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_5_downstream_latency_counter <= p1_std_2s60_burst_5_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_5_downstream_latency_counter = ((std_2s60_burst_5_downstream_run & std_2s60_burst_5_downstream_read))? latency_load_value :
    (std_2s60_burst_5_downstream_latency_counter)? std_2s60_burst_5_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {std_2s60_burst_5_downstream_requests_lan91c111_s1}} & 2) |
    ({2 {std_2s60_burst_5_downstream_requests_ext_ram_s1}} & 2);

  //std_2s60_burst_5_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_5_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_5_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_address_last_time <= std_2s60_burst_5_downstream_address;
    end


  //std_2s60_burst_5/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_5_downstream_waitrequest & (std_2s60_burst_5_downstream_read | std_2s60_burst_5_downstream_write);
    end


  //std_2s60_burst_5_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_address != std_2s60_burst_5_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_5_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_burstcount_last_time <= std_2s60_burst_5_downstream_burstcount;
    end


  //std_2s60_burst_5_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_burstcount != std_2s60_burst_5_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_5_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_byteenable_last_time <= std_2s60_burst_5_downstream_byteenable;
    end


  //std_2s60_burst_5_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_byteenable != std_2s60_burst_5_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_5_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_read_last_time <= std_2s60_burst_5_downstream_read;
    end


  //std_2s60_burst_5_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_read != std_2s60_burst_5_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_5_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_write_last_time <= std_2s60_burst_5_downstream_write;
    end


  //std_2s60_burst_5_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_write != std_2s60_burst_5_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_5_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_5_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_5_downstream_writedata_last_time <= std_2s60_burst_5_downstream_writedata;
    end


  //std_2s60_burst_5_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_5_downstream_writedata != std_2s60_burst_5_downstream_writedata_last_time) & std_2s60_burst_5_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_5_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_6_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_6_upstream_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_6_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_instruction_master_address_to_slave,
                                               cpu_instruction_master_burstcount,
                                               cpu_instruction_master_latency_counter,
                                               cpu_instruction_master_read,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                               reset_n,
                                               std_2s60_burst_6_upstream_readdata,
                                               std_2s60_burst_6_upstream_readdatavalid,
                                               std_2s60_burst_6_upstream_waitrequest,

                                              // outputs:
                                               cpu_instruction_master_granted_std_2s60_burst_6_upstream,
                                               cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                               cpu_instruction_master_requests_std_2s60_burst_6_upstream,
                                               d1_std_2s60_burst_6_upstream_end_xfer,
                                               std_2s60_burst_6_upstream_address,
                                               std_2s60_burst_6_upstream_byteaddress,
                                               std_2s60_burst_6_upstream_byteenable,
                                               std_2s60_burst_6_upstream_debugaccess,
                                               std_2s60_burst_6_upstream_read,
                                               std_2s60_burst_6_upstream_readdata_from_sa,
                                               std_2s60_burst_6_upstream_waitrequest_from_sa,
                                               std_2s60_burst_6_upstream_write
                                            )
;

  output           cpu_instruction_master_granted_std_2s60_burst_6_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_6_upstream;
  output           d1_std_2s60_burst_6_upstream_end_xfer;
  output  [ 15: 0] std_2s60_burst_6_upstream_address;
  output  [ 17: 0] std_2s60_burst_6_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_6_upstream_byteenable;
  output           std_2s60_burst_6_upstream_debugaccess;
  output           std_2s60_burst_6_upstream_read;
  output  [ 31: 0] std_2s60_burst_6_upstream_readdata_from_sa;
  output           std_2s60_burst_6_upstream_waitrequest_from_sa;
  output           std_2s60_burst_6_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_6_upstream_readdata;
  input            std_2s60_burst_6_upstream_readdatavalid;
  input            std_2s60_burst_6_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_6_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_6_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_6_upstream_load_fifo;
  wire    [ 15: 0] std_2s60_burst_6_upstream_address;
  wire             std_2s60_burst_6_upstream_allgrants;
  wire             std_2s60_burst_6_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_6_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_6_upstream_any_continuerequest;
  wire             std_2s60_burst_6_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_6_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_6_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_6_upstream_arb_share_set_values;
  wire             std_2s60_burst_6_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_6_upstream_begins_xfer;
  wire             std_2s60_burst_6_upstream_burstcount_fifo_empty;
  wire    [ 17: 0] std_2s60_burst_6_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_6_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_6_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_6_upstream_current_burst_minus_one;
  wire             std_2s60_burst_6_upstream_debugaccess;
  wire             std_2s60_burst_6_upstream_end_xfer;
  wire             std_2s60_burst_6_upstream_firsttransfer;
  wire             std_2s60_burst_6_upstream_grant_vector;
  wire             std_2s60_burst_6_upstream_in_a_read_cycle;
  wire             std_2s60_burst_6_upstream_in_a_write_cycle;
  reg              std_2s60_burst_6_upstream_load_fifo;
  wire             std_2s60_burst_6_upstream_master_qreq_vector;
  wire             std_2s60_burst_6_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_6_upstream_next_burst_count;
  wire             std_2s60_burst_6_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_6_upstream_read;
  wire    [ 31: 0] std_2s60_burst_6_upstream_readdata_from_sa;
  wire             std_2s60_burst_6_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_6_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_6_upstream_selected_burstcount;
  reg              std_2s60_burst_6_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_6_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_6_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_6_upstream_transaction_burst_count;
  wire             std_2s60_burst_6_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_6_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_6_upstream_waits_for_read;
  wire             std_2s60_burst_6_upstream_waits_for_write;
  wire             std_2s60_burst_6_upstream_write;
  wire             wait_for_std_2s60_burst_6_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_6_upstream_end_xfer;
    end


  assign std_2s60_burst_6_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream));
  //assign std_2s60_burst_6_upstream_readdatavalid_from_sa = std_2s60_burst_6_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_6_upstream_readdatavalid_from_sa = std_2s60_burst_6_upstream_readdatavalid;

  //assign std_2s60_burst_6_upstream_readdata_from_sa = std_2s60_burst_6_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_6_upstream_readdata_from_sa = std_2s60_burst_6_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_6_upstream = (({cpu_instruction_master_address_to_slave[25 : 16] , 16'b0} == 26'h2120000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_6_upstream_waitrequest_from_sa = std_2s60_burst_6_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_6_upstream_waitrequest_from_sa = std_2s60_burst_6_upstream_waitrequest;

  //std_2s60_burst_6_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_6_upstream_arb_share_set_values = 1;

  //std_2s60_burst_6_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_6_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_6_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_6_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_6_upstream;

  //std_2s60_burst_6_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_6_upstream_arb_share_counter_next_value = std_2s60_burst_6_upstream_firsttransfer ? (std_2s60_burst_6_upstream_arb_share_set_values - 1) : |std_2s60_burst_6_upstream_arb_share_counter ? (std_2s60_burst_6_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_6_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_6_upstream_allgrants = |std_2s60_burst_6_upstream_grant_vector;

  //std_2s60_burst_6_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_6_upstream_end_xfer = ~(std_2s60_burst_6_upstream_waits_for_read | std_2s60_burst_6_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream = std_2s60_burst_6_upstream_end_xfer & (~std_2s60_burst_6_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_6_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_6_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream & std_2s60_burst_6_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream & ~std_2s60_burst_6_upstream_non_bursting_master_requests);

  //std_2s60_burst_6_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_6_upstream_arb_counter_enable)
          std_2s60_burst_6_upstream_arb_share_counter <= std_2s60_burst_6_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_6_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_6_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_6_upstream & ~std_2s60_burst_6_upstream_non_bursting_master_requests))
          std_2s60_burst_6_upstream_slavearbiterlockenable <= |std_2s60_burst_6_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_6/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_6_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_6_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_6_upstream_slavearbiterlockenable2 = |std_2s60_burst_6_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_6/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_6_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_6_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_6_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream = cpu_instruction_master_requests_std_2s60_burst_6_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register))));
  //unique name for std_2s60_burst_6_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_6_upstream_move_on_to_next_transaction = std_2s60_burst_6_upstream_this_cycle_is_the_last_burst & std_2s60_burst_6_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_6_upstream, which is an e_mux
  assign std_2s60_burst_6_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_6_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_6_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_6_upstream_module burstcount_fifo_for_std_2s60_burst_6_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_6_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_6_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_6_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_6_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read & std_2s60_burst_6_upstream_load_fifo & ~(std_2s60_burst_6_upstream_this_cycle_is_the_last_burst & std_2s60_burst_6_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_6_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_6_upstream_current_burst_minus_one = std_2s60_burst_6_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_6_upstream, which is an e_mux
  assign std_2s60_burst_6_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read) & ~std_2s60_burst_6_upstream_load_fifo))? std_2s60_burst_6_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read & std_2s60_burst_6_upstream_this_cycle_is_the_last_burst & std_2s60_burst_6_upstream_burstcount_fifo_empty))? std_2s60_burst_6_upstream_selected_burstcount :
    (std_2s60_burst_6_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_6_upstream_transaction_burst_count :
    std_2s60_burst_6_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_6_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_upstream_current_burst <= 0;
      else if (std_2s60_burst_6_upstream_readdatavalid_from_sa | (~std_2s60_burst_6_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read)))
          std_2s60_burst_6_upstream_current_burst <= std_2s60_burst_6_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_6_upstream_load_fifo = (~std_2s60_burst_6_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read) & std_2s60_burst_6_upstream_load_fifo))? 1 :
    ~std_2s60_burst_6_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read) & ~std_2s60_burst_6_upstream_load_fifo | std_2s60_burst_6_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_6_upstream_load_fifo <= p0_std_2s60_burst_6_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_6_upstream, which is an e_assign
  assign std_2s60_burst_6_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_6_upstream_current_burst_minus_one) & std_2s60_burst_6_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_6_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_6_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_6_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_6_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_6_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_6_upstream),
      .full                 (),
      .read                 (std_2s60_burst_6_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_6_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_6_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream = std_2s60_burst_6_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_6/upstream, which is an e_mux
  assign std_2s60_burst_6_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_6_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_6/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_6_upstream = cpu_instruction_master_requests_std_2s60_burst_6_upstream;

  //allow new arb cycle for std_2s60_burst_6/upstream, which is an e_assign
  assign std_2s60_burst_6_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_6_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_6_upstream_master_qreq_vector = 1;

  //std_2s60_burst_6_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_6_upstream_firsttransfer = std_2s60_burst_6_upstream_begins_xfer ? std_2s60_burst_6_upstream_unreg_firsttransfer : std_2s60_burst_6_upstream_reg_firsttransfer;

  //std_2s60_burst_6_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_6_upstream_unreg_firsttransfer = ~(std_2s60_burst_6_upstream_slavearbiterlockenable & std_2s60_burst_6_upstream_any_continuerequest);

  //std_2s60_burst_6_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_6_upstream_begins_xfer)
          std_2s60_burst_6_upstream_reg_firsttransfer <= std_2s60_burst_6_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_6_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_6_upstream_beginbursttransfer_internal = std_2s60_burst_6_upstream_begins_xfer;

  //std_2s60_burst_6_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_6_upstream_read = cpu_instruction_master_granted_std_2s60_burst_6_upstream & cpu_instruction_master_read;

  //std_2s60_burst_6_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_6_upstream_write = 0;

  //std_2s60_burst_6_upstream_address mux, which is an e_mux
  assign std_2s60_burst_6_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_std_2s60_burst_6_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_6_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_6_upstream_end_xfer <= std_2s60_burst_6_upstream_end_xfer;
    end


  //std_2s60_burst_6_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_6_upstream_waits_for_read = std_2s60_burst_6_upstream_in_a_read_cycle & std_2s60_burst_6_upstream_waitrequest_from_sa;

  //std_2s60_burst_6_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_6_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_6_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_6_upstream_in_a_read_cycle;

  //std_2s60_burst_6_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_6_upstream_waits_for_write = std_2s60_burst_6_upstream_in_a_write_cycle & std_2s60_burst_6_upstream_waitrequest_from_sa;

  //std_2s60_burst_6_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_6_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_6_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_6_upstream_counter = 0;
  //std_2s60_burst_6_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_6_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_6_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_6/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_6_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_6/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_6_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_onchip_ram_64_kbytes_s1_end_xfer,
                                                 onchip_ram_64_kbytes_s1_readdata_from_sa,
                                                 reset_n,
                                                 std_2s60_burst_6_downstream_address,
                                                 std_2s60_burst_6_downstream_burstcount,
                                                 std_2s60_burst_6_downstream_byteenable,
                                                 std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_6_downstream_read,
                                                 std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_6_downstream_write,
                                                 std_2s60_burst_6_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_6_downstream_address_to_slave,
                                                 std_2s60_burst_6_downstream_latency_counter,
                                                 std_2s60_burst_6_downstream_readdata,
                                                 std_2s60_burst_6_downstream_readdatavalid,
                                                 std_2s60_burst_6_downstream_reset_n,
                                                 std_2s60_burst_6_downstream_waitrequest
                                              )
;

  output  [ 15: 0] std_2s60_burst_6_downstream_address_to_slave;
  output           std_2s60_burst_6_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_6_downstream_readdata;
  output           std_2s60_burst_6_downstream_readdatavalid;
  output           std_2s60_burst_6_downstream_reset_n;
  output           std_2s60_burst_6_downstream_waitrequest;
  input            clk;
  input            d1_onchip_ram_64_kbytes_s1_end_xfer;
  input   [ 31: 0] onchip_ram_64_kbytes_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_6_downstream_address;
  input            std_2s60_burst_6_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_6_downstream_byteenable;
  input            std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_6_downstream_read;
  input            std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_6_downstream_write;
  input   [ 31: 0] std_2s60_burst_6_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_6_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_6_downstream_readdatavalid;
  wire             r_0;
  reg     [ 15: 0] std_2s60_burst_6_downstream_address_last_time;
  wire    [ 15: 0] std_2s60_burst_6_downstream_address_to_slave;
  reg              std_2s60_burst_6_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_6_downstream_byteenable_last_time;
  wire             std_2s60_burst_6_downstream_is_granted_some_slave;
  reg              std_2s60_burst_6_downstream_latency_counter;
  reg              std_2s60_burst_6_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_6_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_6_downstream_readdata;
  wire             std_2s60_burst_6_downstream_readdatavalid;
  wire             std_2s60_burst_6_downstream_reset_n;
  wire             std_2s60_burst_6_downstream_run;
  wire             std_2s60_burst_6_downstream_waitrequest;
  reg              std_2s60_burst_6_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_6_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1) & (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1 | ~std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1) & ((~std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~(std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write) | (1 & (std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write)))) & ((~std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~(std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write) | (1 & (std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_6_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_6_downstream_address_to_slave = std_2s60_burst_6_downstream_address;

  //std_2s60_burst_6_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_6_downstream_read_but_no_slave_selected <= std_2s60_burst_6_downstream_read & std_2s60_burst_6_downstream_run & ~std_2s60_burst_6_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_6_downstream_is_granted_some_slave = std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_6_downstream_readdatavalid = std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_6_downstream_readdatavalid = std_2s60_burst_6_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_6_downstream_readdatavalid;

  //std_2s60_burst_6/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_6_downstream_readdata = onchip_ram_64_kbytes_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_6_downstream_waitrequest = ~std_2s60_burst_6_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_6_downstream_latency_counter <= p1_std_2s60_burst_6_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_6_downstream_latency_counter = ((std_2s60_burst_6_downstream_run & std_2s60_burst_6_downstream_read))? latency_load_value :
    (std_2s60_burst_6_downstream_latency_counter)? std_2s60_burst_6_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1}} & 1;

  //std_2s60_burst_6_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_6_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_6_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_address_last_time <= std_2s60_burst_6_downstream_address;
    end


  //std_2s60_burst_6/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_6_downstream_waitrequest & (std_2s60_burst_6_downstream_read | std_2s60_burst_6_downstream_write);
    end


  //std_2s60_burst_6_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_address != std_2s60_burst_6_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_6_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_burstcount_last_time <= std_2s60_burst_6_downstream_burstcount;
    end


  //std_2s60_burst_6_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_burstcount != std_2s60_burst_6_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_6_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_byteenable_last_time <= std_2s60_burst_6_downstream_byteenable;
    end


  //std_2s60_burst_6_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_byteenable != std_2s60_burst_6_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_6_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_read_last_time <= std_2s60_burst_6_downstream_read;
    end


  //std_2s60_burst_6_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_read != std_2s60_burst_6_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_6_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_write_last_time <= std_2s60_burst_6_downstream_write;
    end


  //std_2s60_burst_6_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_write != std_2s60_burst_6_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_6_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_6_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_6_downstream_writedata_last_time <= std_2s60_burst_6_downstream_writedata;
    end


  //std_2s60_burst_6_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_6_downstream_writedata != std_2s60_burst_6_downstream_writedata_last_time) & std_2s60_burst_6_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_6_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_7_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_7_upstream_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_7_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_burstcount,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_debugaccess,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                               cpu_data_master_write,
                                               cpu_data_master_writedata,
                                               reset_n,
                                               std_2s60_burst_7_upstream_readdata,
                                               std_2s60_burst_7_upstream_readdatavalid,
                                               std_2s60_burst_7_upstream_waitrequest,

                                              // outputs:
                                               cpu_data_master_granted_std_2s60_burst_7_upstream,
                                               cpu_data_master_qualified_request_std_2s60_burst_7_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                               cpu_data_master_requests_std_2s60_burst_7_upstream,
                                               d1_std_2s60_burst_7_upstream_end_xfer,
                                               std_2s60_burst_7_upstream_address,
                                               std_2s60_burst_7_upstream_burstcount,
                                               std_2s60_burst_7_upstream_byteaddress,
                                               std_2s60_burst_7_upstream_byteenable,
                                               std_2s60_burst_7_upstream_debugaccess,
                                               std_2s60_burst_7_upstream_read,
                                               std_2s60_burst_7_upstream_readdata_from_sa,
                                               std_2s60_burst_7_upstream_waitrequest_from_sa,
                                               std_2s60_burst_7_upstream_write,
                                               std_2s60_burst_7_upstream_writedata
                                            )
;

  output           cpu_data_master_granted_std_2s60_burst_7_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_7_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_7_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_7_upstream;
  output           d1_std_2s60_burst_7_upstream_end_xfer;
  output  [ 15: 0] std_2s60_burst_7_upstream_address;
  output  [  3: 0] std_2s60_burst_7_upstream_burstcount;
  output  [ 17: 0] std_2s60_burst_7_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_7_upstream_byteenable;
  output           std_2s60_burst_7_upstream_debugaccess;
  output           std_2s60_burst_7_upstream_read;
  output  [ 31: 0] std_2s60_burst_7_upstream_readdata_from_sa;
  output           std_2s60_burst_7_upstream_waitrequest_from_sa;
  output           std_2s60_burst_7_upstream_write;
  output  [ 31: 0] std_2s60_burst_7_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_7_upstream_readdata;
  input            std_2s60_burst_7_upstream_readdatavalid;
  input            std_2s60_burst_7_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_7_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_7_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_7_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_7_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_7_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_7_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_7_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_7_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_7_upstream_load_fifo;
  wire    [ 15: 0] std_2s60_burst_7_upstream_address;
  wire             std_2s60_burst_7_upstream_allgrants;
  wire             std_2s60_burst_7_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_7_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_7_upstream_any_continuerequest;
  wire             std_2s60_burst_7_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_7_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_7_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_7_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_7_upstream_bbt_burstcounter;
  wire             std_2s60_burst_7_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_7_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_7_upstream_burstcount;
  wire             std_2s60_burst_7_upstream_burstcount_fifo_empty;
  wire    [ 17: 0] std_2s60_burst_7_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_7_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_7_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_7_upstream_current_burst_minus_one;
  wire             std_2s60_burst_7_upstream_debugaccess;
  wire             std_2s60_burst_7_upstream_end_xfer;
  wire             std_2s60_burst_7_upstream_firsttransfer;
  wire             std_2s60_burst_7_upstream_grant_vector;
  wire             std_2s60_burst_7_upstream_in_a_read_cycle;
  wire             std_2s60_burst_7_upstream_in_a_write_cycle;
  reg              std_2s60_burst_7_upstream_load_fifo;
  wire             std_2s60_burst_7_upstream_master_qreq_vector;
  wire             std_2s60_burst_7_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_7_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_7_upstream_next_burst_count;
  wire             std_2s60_burst_7_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_7_upstream_read;
  wire    [ 31: 0] std_2s60_burst_7_upstream_readdata_from_sa;
  wire             std_2s60_burst_7_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_7_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_7_upstream_selected_burstcount;
  reg              std_2s60_burst_7_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_7_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_7_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_7_upstream_transaction_burst_count;
  wire             std_2s60_burst_7_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_7_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_7_upstream_waits_for_read;
  wire             std_2s60_burst_7_upstream_waits_for_write;
  wire             std_2s60_burst_7_upstream_write;
  wire    [ 31: 0] std_2s60_burst_7_upstream_writedata;
  wire             wait_for_std_2s60_burst_7_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_7_upstream_end_xfer;
    end


  assign std_2s60_burst_7_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_7_upstream));
  //assign std_2s60_burst_7_upstream_readdatavalid_from_sa = std_2s60_burst_7_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_7_upstream_readdatavalid_from_sa = std_2s60_burst_7_upstream_readdatavalid;

  //assign std_2s60_burst_7_upstream_readdata_from_sa = std_2s60_burst_7_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_7_upstream_readdata_from_sa = std_2s60_burst_7_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_7_upstream = ({cpu_data_master_address_to_slave[25 : 16] , 16'b0} == 26'h2120000) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_7_upstream_waitrequest_from_sa = std_2s60_burst_7_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_7_upstream_waitrequest_from_sa = std_2s60_burst_7_upstream_waitrequest;

  //std_2s60_burst_7_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_7_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_7_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_7_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_7_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_7_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_7_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_7_upstream;

  //std_2s60_burst_7_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_7_upstream_arb_share_counter_next_value = std_2s60_burst_7_upstream_firsttransfer ? (std_2s60_burst_7_upstream_arb_share_set_values - 1) : |std_2s60_burst_7_upstream_arb_share_counter ? (std_2s60_burst_7_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_7_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_7_upstream_allgrants = |std_2s60_burst_7_upstream_grant_vector;

  //std_2s60_burst_7_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_7_upstream_end_xfer = ~(std_2s60_burst_7_upstream_waits_for_read | std_2s60_burst_7_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream = std_2s60_burst_7_upstream_end_xfer & (~std_2s60_burst_7_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_7_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_7_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream & std_2s60_burst_7_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream & ~std_2s60_burst_7_upstream_non_bursting_master_requests);

  //std_2s60_burst_7_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_7_upstream_arb_counter_enable)
          std_2s60_burst_7_upstream_arb_share_counter <= std_2s60_burst_7_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_7_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_7_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_7_upstream & ~std_2s60_burst_7_upstream_non_bursting_master_requests))
          std_2s60_burst_7_upstream_slavearbiterlockenable <= |std_2s60_burst_7_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_7/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_7_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_7_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_7_upstream_slavearbiterlockenable2 = |std_2s60_burst_7_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_7/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_7_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_7_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_7_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_7_upstream = cpu_data_master_requests_std_2s60_burst_7_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register))));
  //unique name for std_2s60_burst_7_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_7_upstream_move_on_to_next_transaction = std_2s60_burst_7_upstream_this_cycle_is_the_last_burst & std_2s60_burst_7_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_7_upstream, which is an e_mux
  assign std_2s60_burst_7_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_7_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_7_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_7_upstream_module burstcount_fifo_for_std_2s60_burst_7_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_7_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_7_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_7_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_7_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read & std_2s60_burst_7_upstream_load_fifo & ~(std_2s60_burst_7_upstream_this_cycle_is_the_last_burst & std_2s60_burst_7_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_7_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_7_upstream_current_burst_minus_one = std_2s60_burst_7_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_7_upstream, which is an e_mux
  assign std_2s60_burst_7_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read) & ~std_2s60_burst_7_upstream_load_fifo))? std_2s60_burst_7_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read & std_2s60_burst_7_upstream_this_cycle_is_the_last_burst & std_2s60_burst_7_upstream_burstcount_fifo_empty))? std_2s60_burst_7_upstream_selected_burstcount :
    (std_2s60_burst_7_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_7_upstream_transaction_burst_count :
    std_2s60_burst_7_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_7_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_current_burst <= 0;
      else if (std_2s60_burst_7_upstream_readdatavalid_from_sa | (~std_2s60_burst_7_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read)))
          std_2s60_burst_7_upstream_current_burst <= std_2s60_burst_7_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_7_upstream_load_fifo = (~std_2s60_burst_7_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read) & std_2s60_burst_7_upstream_load_fifo))? 1 :
    ~std_2s60_burst_7_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read) & ~std_2s60_burst_7_upstream_load_fifo | std_2s60_burst_7_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_7_upstream_load_fifo <= p0_std_2s60_burst_7_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_7_upstream, which is an e_assign
  assign std_2s60_burst_7_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_7_upstream_current_burst_minus_one) & std_2s60_burst_7_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_7_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_7_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_7_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_7_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_7_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_7_upstream),
      .full                 (),
      .read                 (std_2s60_burst_7_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_7_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_7_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_7_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_7_upstream = std_2s60_burst_7_upstream_readdatavalid_from_sa;

  //std_2s60_burst_7_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_7_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_7/upstream, which is an e_mux
  assign std_2s60_burst_7_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_7_upstream = cpu_data_master_qualified_request_std_2s60_burst_7_upstream;

  //cpu/data_master saved-grant std_2s60_burst_7/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_7_upstream = cpu_data_master_requests_std_2s60_burst_7_upstream;

  //allow new arb cycle for std_2s60_burst_7/upstream, which is an e_assign
  assign std_2s60_burst_7_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_7_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_7_upstream_master_qreq_vector = 1;

  //std_2s60_burst_7_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_7_upstream_firsttransfer = std_2s60_burst_7_upstream_begins_xfer ? std_2s60_burst_7_upstream_unreg_firsttransfer : std_2s60_burst_7_upstream_reg_firsttransfer;

  //std_2s60_burst_7_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_7_upstream_unreg_firsttransfer = ~(std_2s60_burst_7_upstream_slavearbiterlockenable & std_2s60_burst_7_upstream_any_continuerequest);

  //std_2s60_burst_7_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_7_upstream_begins_xfer)
          std_2s60_burst_7_upstream_reg_firsttransfer <= std_2s60_burst_7_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_7_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_7_upstream_next_bbt_burstcount = ((((std_2s60_burst_7_upstream_write) && (std_2s60_burst_7_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_7_upstream_burstcount - 1) :
    ((((std_2s60_burst_7_upstream_read) && (std_2s60_burst_7_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_7_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_7_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_7_upstream_begins_xfer)
          std_2s60_burst_7_upstream_bbt_burstcounter <= std_2s60_burst_7_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_7_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_7_upstream_beginbursttransfer_internal = std_2s60_burst_7_upstream_begins_xfer & (std_2s60_burst_7_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_7_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_7_upstream_read = cpu_data_master_granted_std_2s60_burst_7_upstream & cpu_data_master_read;

  //std_2s60_burst_7_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_7_upstream_write = cpu_data_master_granted_std_2s60_burst_7_upstream & cpu_data_master_write;

  //std_2s60_burst_7_upstream_address mux, which is an e_mux
  assign std_2s60_burst_7_upstream_address = cpu_data_master_address_to_slave;

  //d1_std_2s60_burst_7_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_7_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_7_upstream_end_xfer <= std_2s60_burst_7_upstream_end_xfer;
    end


  //std_2s60_burst_7_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_7_upstream_waits_for_read = std_2s60_burst_7_upstream_in_a_read_cycle & std_2s60_burst_7_upstream_waitrequest_from_sa;

  //std_2s60_burst_7_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_7_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_7_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_7_upstream_in_a_read_cycle;

  //std_2s60_burst_7_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_7_upstream_waits_for_write = std_2s60_burst_7_upstream_in_a_write_cycle & std_2s60_burst_7_upstream_waitrequest_from_sa;

  //std_2s60_burst_7_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_7_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_7_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_7_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_7_upstream_counter = 0;
  //std_2s60_burst_7_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_7_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_7_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_7_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_7_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_7_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_7_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_7/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_7_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_7/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_7_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_onchip_ram_64_kbytes_s1_end_xfer,
                                                 onchip_ram_64_kbytes_s1_readdata_from_sa,
                                                 reset_n,
                                                 std_2s60_burst_7_downstream_address,
                                                 std_2s60_burst_7_downstream_burstcount,
                                                 std_2s60_burst_7_downstream_byteenable,
                                                 std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_7_downstream_read,
                                                 std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1,
                                                 std_2s60_burst_7_downstream_write,
                                                 std_2s60_burst_7_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_7_downstream_address_to_slave,
                                                 std_2s60_burst_7_downstream_latency_counter,
                                                 std_2s60_burst_7_downstream_readdata,
                                                 std_2s60_burst_7_downstream_readdatavalid,
                                                 std_2s60_burst_7_downstream_reset_n,
                                                 std_2s60_burst_7_downstream_waitrequest
                                              )
;

  output  [ 15: 0] std_2s60_burst_7_downstream_address_to_slave;
  output           std_2s60_burst_7_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_7_downstream_readdata;
  output           std_2s60_burst_7_downstream_readdatavalid;
  output           std_2s60_burst_7_downstream_reset_n;
  output           std_2s60_burst_7_downstream_waitrequest;
  input            clk;
  input            d1_onchip_ram_64_kbytes_s1_end_xfer;
  input   [ 31: 0] onchip_ram_64_kbytes_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_7_downstream_address;
  input            std_2s60_burst_7_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_7_downstream_byteenable;
  input            std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_7_downstream_read;
  input            std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1;
  input            std_2s60_burst_7_downstream_write;
  input   [ 31: 0] std_2s60_burst_7_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_std_2s60_burst_7_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_7_downstream_readdatavalid;
  wire             r_0;
  reg     [ 15: 0] std_2s60_burst_7_downstream_address_last_time;
  wire    [ 15: 0] std_2s60_burst_7_downstream_address_to_slave;
  reg              std_2s60_burst_7_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_7_downstream_byteenable_last_time;
  wire             std_2s60_burst_7_downstream_is_granted_some_slave;
  reg              std_2s60_burst_7_downstream_latency_counter;
  reg              std_2s60_burst_7_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_7_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_7_downstream_readdata;
  wire             std_2s60_burst_7_downstream_readdatavalid;
  wire             std_2s60_burst_7_downstream_reset_n;
  wire             std_2s60_burst_7_downstream_run;
  wire             std_2s60_burst_7_downstream_waitrequest;
  reg              std_2s60_burst_7_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_7_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1) & (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1 | ~std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1) & ((~std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~(std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write) | (1 & (std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write)))) & ((~std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 | ~(std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write) | (1 & (std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_7_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_7_downstream_address_to_slave = std_2s60_burst_7_downstream_address;

  //std_2s60_burst_7_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_7_downstream_read_but_no_slave_selected <= std_2s60_burst_7_downstream_read & std_2s60_burst_7_downstream_run & ~std_2s60_burst_7_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_7_downstream_is_granted_some_slave = std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_7_downstream_readdatavalid = std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_7_downstream_readdatavalid = std_2s60_burst_7_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_7_downstream_readdatavalid;

  //std_2s60_burst_7/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_7_downstream_readdata = onchip_ram_64_kbytes_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_7_downstream_waitrequest = ~std_2s60_burst_7_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_7_downstream_latency_counter <= p1_std_2s60_burst_7_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_7_downstream_latency_counter = ((std_2s60_burst_7_downstream_run & std_2s60_burst_7_downstream_read))? latency_load_value :
    (std_2s60_burst_7_downstream_latency_counter)? std_2s60_burst_7_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1}} & 1;

  //std_2s60_burst_7_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_7_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_7_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_address_last_time <= std_2s60_burst_7_downstream_address;
    end


  //std_2s60_burst_7/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_7_downstream_waitrequest & (std_2s60_burst_7_downstream_read | std_2s60_burst_7_downstream_write);
    end


  //std_2s60_burst_7_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_address != std_2s60_burst_7_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_7_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_burstcount_last_time <= std_2s60_burst_7_downstream_burstcount;
    end


  //std_2s60_burst_7_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_burstcount != std_2s60_burst_7_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_7_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_byteenable_last_time <= std_2s60_burst_7_downstream_byteenable;
    end


  //std_2s60_burst_7_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_byteenable != std_2s60_burst_7_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_7_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_read_last_time <= std_2s60_burst_7_downstream_read;
    end


  //std_2s60_burst_7_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_read != std_2s60_burst_7_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_7_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_write_last_time <= std_2s60_burst_7_downstream_write;
    end


  //std_2s60_burst_7_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_write != std_2s60_burst_7_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_7_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_7_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_7_downstream_writedata_last_time <= std_2s60_burst_7_downstream_writedata;
    end


  //std_2s60_burst_7_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_7_downstream_writedata != std_2s60_burst_7_downstream_writedata_last_time) & std_2s60_burst_7_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_7_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_8_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_8_upstream_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_8_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_instruction_master_address_to_slave,
                                               cpu_instruction_master_burstcount,
                                               cpu_instruction_master_latency_counter,
                                               cpu_instruction_master_read,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register,
                                               reset_n,
                                               std_2s60_burst_8_upstream_readdata,
                                               std_2s60_burst_8_upstream_readdatavalid,
                                               std_2s60_burst_8_upstream_waitrequest,

                                              // outputs:
                                               cpu_instruction_master_granted_std_2s60_burst_8_upstream,
                                               cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream,
                                               cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register,
                                               cpu_instruction_master_requests_std_2s60_burst_8_upstream,
                                               d1_std_2s60_burst_8_upstream_end_xfer,
                                               std_2s60_burst_8_upstream_address,
                                               std_2s60_burst_8_upstream_byteaddress,
                                               std_2s60_burst_8_upstream_byteenable,
                                               std_2s60_burst_8_upstream_debugaccess,
                                               std_2s60_burst_8_upstream_read,
                                               std_2s60_burst_8_upstream_readdata_from_sa,
                                               std_2s60_burst_8_upstream_waitrequest_from_sa,
                                               std_2s60_burst_8_upstream_write
                                            )
;

  output           cpu_instruction_master_granted_std_2s60_burst_8_upstream;
  output           cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream;
  output           cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  output           cpu_instruction_master_requests_std_2s60_burst_8_upstream;
  output           d1_std_2s60_burst_8_upstream_end_xfer;
  output  [ 15: 0] std_2s60_burst_8_upstream_address;
  output  [ 17: 0] std_2s60_burst_8_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_8_upstream_byteenable;
  output           std_2s60_burst_8_upstream_debugaccess;
  output           std_2s60_burst_8_upstream_read;
  output  [ 31: 0] std_2s60_burst_8_upstream_readdata_from_sa;
  output           std_2s60_burst_8_upstream_waitrequest_from_sa;
  output           std_2s60_burst_8_upstream_write;
  input            clk;
  input   [ 25: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_8_upstream_readdata;
  input            std_2s60_burst_8_upstream_readdatavalid;
  input            std_2s60_burst_8_upstream_waitrequest;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  wire             cpu_instruction_master_requests_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_saved_grant_std_2s60_burst_8_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_8_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_8_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_8_upstream_from_cpu_instruction_master;
  wire    [ 15: 0] std_2s60_burst_8_upstream_address;
  wire             std_2s60_burst_8_upstream_allgrants;
  wire             std_2s60_burst_8_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_8_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_8_upstream_any_continuerequest;
  wire             std_2s60_burst_8_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_8_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_8_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_8_upstream_arb_share_set_values;
  wire             std_2s60_burst_8_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_8_upstream_begins_xfer;
  wire             std_2s60_burst_8_upstream_burstcount_fifo_empty;
  wire    [ 17: 0] std_2s60_burst_8_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_8_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_8_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_8_upstream_current_burst_minus_one;
  wire             std_2s60_burst_8_upstream_debugaccess;
  wire             std_2s60_burst_8_upstream_end_xfer;
  wire             std_2s60_burst_8_upstream_firsttransfer;
  wire             std_2s60_burst_8_upstream_grant_vector;
  wire             std_2s60_burst_8_upstream_in_a_read_cycle;
  wire             std_2s60_burst_8_upstream_in_a_write_cycle;
  reg              std_2s60_burst_8_upstream_load_fifo;
  wire             std_2s60_burst_8_upstream_master_qreq_vector;
  wire             std_2s60_burst_8_upstream_move_on_to_next_transaction;
  wire    [  3: 0] std_2s60_burst_8_upstream_next_burst_count;
  wire             std_2s60_burst_8_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_8_upstream_read;
  wire    [ 31: 0] std_2s60_burst_8_upstream_readdata_from_sa;
  wire             std_2s60_burst_8_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_8_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_8_upstream_selected_burstcount;
  reg              std_2s60_burst_8_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_8_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_8_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_8_upstream_transaction_burst_count;
  wire             std_2s60_burst_8_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_8_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_8_upstream_waits_for_read;
  wire             std_2s60_burst_8_upstream_waits_for_write;
  wire             std_2s60_burst_8_upstream_write;
  wire             wait_for_std_2s60_burst_8_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_8_upstream_end_xfer;
    end


  assign std_2s60_burst_8_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream));
  //assign std_2s60_burst_8_upstream_readdatavalid_from_sa = std_2s60_burst_8_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_8_upstream_readdatavalid_from_sa = std_2s60_burst_8_upstream_readdatavalid;

  //assign std_2s60_burst_8_upstream_readdata_from_sa = std_2s60_burst_8_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_8_upstream_readdata_from_sa = std_2s60_burst_8_upstream_readdata;

  assign cpu_instruction_master_requests_std_2s60_burst_8_upstream = (({cpu_instruction_master_address_to_slave[25 : 16] , 16'b0} == 26'h2110000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign std_2s60_burst_8_upstream_waitrequest_from_sa = std_2s60_burst_8_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_8_upstream_waitrequest_from_sa = std_2s60_burst_8_upstream_waitrequest;

  //std_2s60_burst_8_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_8_upstream_arb_share_set_values = 1;

  //std_2s60_burst_8_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_8_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_8_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_8_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_std_2s60_burst_8_upstream;

  //std_2s60_burst_8_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_8_upstream_arb_share_counter_next_value = std_2s60_burst_8_upstream_firsttransfer ? (std_2s60_burst_8_upstream_arb_share_set_values - 1) : |std_2s60_burst_8_upstream_arb_share_counter ? (std_2s60_burst_8_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_8_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_8_upstream_allgrants = |std_2s60_burst_8_upstream_grant_vector;

  //std_2s60_burst_8_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_8_upstream_end_xfer = ~(std_2s60_burst_8_upstream_waits_for_read | std_2s60_burst_8_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream = std_2s60_burst_8_upstream_end_xfer & (~std_2s60_burst_8_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_8_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_8_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream & std_2s60_burst_8_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream & ~std_2s60_burst_8_upstream_non_bursting_master_requests);

  //std_2s60_burst_8_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_8_upstream_arb_counter_enable)
          std_2s60_burst_8_upstream_arb_share_counter <= std_2s60_burst_8_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_8_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_8_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_8_upstream & ~std_2s60_burst_8_upstream_non_bursting_master_requests))
          std_2s60_burst_8_upstream_slavearbiterlockenable <= |std_2s60_burst_8_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master std_2s60_burst_8/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = std_2s60_burst_8_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //std_2s60_burst_8_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_8_upstream_slavearbiterlockenable2 = |std_2s60_burst_8_upstream_arb_share_counter_next_value;

  //cpu/instruction_master std_2s60_burst_8/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = std_2s60_burst_8_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //std_2s60_burst_8_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_8_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream = cpu_instruction_master_requests_std_2s60_burst_8_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register) | (|cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register))));
  //unique name for std_2s60_burst_8_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_8_upstream_move_on_to_next_transaction = std_2s60_burst_8_upstream_this_cycle_is_the_last_burst & std_2s60_burst_8_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_8_upstream, which is an e_mux
  assign std_2s60_burst_8_upstream_selected_burstcount = (cpu_instruction_master_granted_std_2s60_burst_8_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_8_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_8_upstream_module burstcount_fifo_for_std_2s60_burst_8_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_8_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_8_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_8_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_8_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read & std_2s60_burst_8_upstream_load_fifo & ~(std_2s60_burst_8_upstream_this_cycle_is_the_last_burst & std_2s60_burst_8_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_8_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_8_upstream_current_burst_minus_one = std_2s60_burst_8_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_8_upstream, which is an e_mux
  assign std_2s60_burst_8_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read) & ~std_2s60_burst_8_upstream_load_fifo))? std_2s60_burst_8_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read & std_2s60_burst_8_upstream_this_cycle_is_the_last_burst & std_2s60_burst_8_upstream_burstcount_fifo_empty))? std_2s60_burst_8_upstream_selected_burstcount :
    (std_2s60_burst_8_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_8_upstream_transaction_burst_count :
    std_2s60_burst_8_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_8_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_upstream_current_burst <= 0;
      else if (std_2s60_burst_8_upstream_readdatavalid_from_sa | (~std_2s60_burst_8_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read)))
          std_2s60_burst_8_upstream_current_burst <= std_2s60_burst_8_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_8_upstream_load_fifo = (~std_2s60_burst_8_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read) & std_2s60_burst_8_upstream_load_fifo))? 1 :
    ~std_2s60_burst_8_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read) & ~std_2s60_burst_8_upstream_load_fifo | std_2s60_burst_8_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_8_upstream_load_fifo <= p0_std_2s60_burst_8_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_8_upstream, which is an e_assign
  assign std_2s60_burst_8_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_8_upstream_current_burst_minus_one) & std_2s60_burst_8_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_8_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_8_upstream_module rdv_fifo_for_cpu_instruction_master_to_std_2s60_burst_8_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_std_2s60_burst_8_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_std_2s60_burst_8_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_8_upstream),
      .full                 (),
      .read                 (std_2s60_burst_8_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_8_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_std_2s60_burst_8_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream = std_2s60_burst_8_upstream_readdatavalid_from_sa;

  //byteaddress mux for std_2s60_burst_8/upstream, which is an e_mux
  assign std_2s60_burst_8_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_std_2s60_burst_8_upstream = cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream;

  //cpu/instruction_master saved-grant std_2s60_burst_8/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_std_2s60_burst_8_upstream = cpu_instruction_master_requests_std_2s60_burst_8_upstream;

  //allow new arb cycle for std_2s60_burst_8/upstream, which is an e_assign
  assign std_2s60_burst_8_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_8_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_8_upstream_master_qreq_vector = 1;

  //std_2s60_burst_8_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_8_upstream_firsttransfer = std_2s60_burst_8_upstream_begins_xfer ? std_2s60_burst_8_upstream_unreg_firsttransfer : std_2s60_burst_8_upstream_reg_firsttransfer;

  //std_2s60_burst_8_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_8_upstream_unreg_firsttransfer = ~(std_2s60_burst_8_upstream_slavearbiterlockenable & std_2s60_burst_8_upstream_any_continuerequest);

  //std_2s60_burst_8_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_8_upstream_begins_xfer)
          std_2s60_burst_8_upstream_reg_firsttransfer <= std_2s60_burst_8_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_8_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_8_upstream_beginbursttransfer_internal = std_2s60_burst_8_upstream_begins_xfer;

  //std_2s60_burst_8_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_8_upstream_read = cpu_instruction_master_granted_std_2s60_burst_8_upstream & cpu_instruction_master_read;

  //std_2s60_burst_8_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_8_upstream_write = 0;

  assign shifted_address_to_std_2s60_burst_8_upstream_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //std_2s60_burst_8_upstream_address mux, which is an e_mux
  assign std_2s60_burst_8_upstream_address = shifted_address_to_std_2s60_burst_8_upstream_from_cpu_instruction_master >> 2;

  //d1_std_2s60_burst_8_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_8_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_8_upstream_end_xfer <= std_2s60_burst_8_upstream_end_xfer;
    end


  //std_2s60_burst_8_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_8_upstream_waits_for_read = std_2s60_burst_8_upstream_in_a_read_cycle & std_2s60_burst_8_upstream_waitrequest_from_sa;

  //std_2s60_burst_8_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_8_upstream_in_a_read_cycle = cpu_instruction_master_granted_std_2s60_burst_8_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_8_upstream_in_a_read_cycle;

  //std_2s60_burst_8_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_8_upstream_waits_for_write = std_2s60_burst_8_upstream_in_a_write_cycle & std_2s60_burst_8_upstream_waitrequest_from_sa;

  //std_2s60_burst_8_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_8_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_8_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_8_upstream_counter = 0;
  //std_2s60_burst_8_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_8_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_8_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_8/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_std_2s60_burst_8_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_8/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_8_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_ram_bus_avalon_slave_end_xfer,
                                                 ext_ram_s1_wait_counter_eq_0,
                                                 incoming_ext_ram_bus_data,
                                                 lan91c111_s1_wait_counter_eq_0,
                                                 reset_n,
                                                 std_2s60_burst_8_downstream_address,
                                                 std_2s60_burst_8_downstream_burstcount,
                                                 std_2s60_burst_8_downstream_byteenable,
                                                 std_2s60_burst_8_downstream_granted_ext_ram_s1,
                                                 std_2s60_burst_8_downstream_granted_lan91c111_s1,
                                                 std_2s60_burst_8_downstream_qualified_request_ext_ram_s1,
                                                 std_2s60_burst_8_downstream_qualified_request_lan91c111_s1,
                                                 std_2s60_burst_8_downstream_read,
                                                 std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1,
                                                 std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1,
                                                 std_2s60_burst_8_downstream_requests_ext_ram_s1,
                                                 std_2s60_burst_8_downstream_requests_lan91c111_s1,
                                                 std_2s60_burst_8_downstream_write,
                                                 std_2s60_burst_8_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_8_downstream_address_to_slave,
                                                 std_2s60_burst_8_downstream_latency_counter,
                                                 std_2s60_burst_8_downstream_readdata,
                                                 std_2s60_burst_8_downstream_readdatavalid,
                                                 std_2s60_burst_8_downstream_reset_n,
                                                 std_2s60_burst_8_downstream_waitrequest
                                              )
;

  output  [ 15: 0] std_2s60_burst_8_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_8_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_8_downstream_readdata;
  output           std_2s60_burst_8_downstream_readdatavalid;
  output           std_2s60_burst_8_downstream_reset_n;
  output           std_2s60_burst_8_downstream_waitrequest;
  input            clk;
  input            d1_ext_ram_bus_avalon_slave_end_xfer;
  input            ext_ram_s1_wait_counter_eq_0;
  input   [ 31: 0] incoming_ext_ram_bus_data;
  input            lan91c111_s1_wait_counter_eq_0;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_8_downstream_address;
  input            std_2s60_burst_8_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_8_downstream_byteenable;
  input            std_2s60_burst_8_downstream_granted_ext_ram_s1;
  input            std_2s60_burst_8_downstream_granted_lan91c111_s1;
  input            std_2s60_burst_8_downstream_qualified_request_ext_ram_s1;
  input            std_2s60_burst_8_downstream_qualified_request_lan91c111_s1;
  input            std_2s60_burst_8_downstream_read;
  input            std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1;
  input            std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1;
  input            std_2s60_burst_8_downstream_requests_ext_ram_s1;
  input            std_2s60_burst_8_downstream_requests_lan91c111_s1;
  input            std_2s60_burst_8_downstream_write;
  input   [ 31: 0] std_2s60_burst_8_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_8_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_8_downstream_readdatavalid;
  wire             r_0;
  reg     [ 15: 0] std_2s60_burst_8_downstream_address_last_time;
  wire    [ 15: 0] std_2s60_burst_8_downstream_address_to_slave;
  reg              std_2s60_burst_8_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_8_downstream_byteenable_last_time;
  wire             std_2s60_burst_8_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_8_downstream_latency_counter;
  reg              std_2s60_burst_8_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_8_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_8_downstream_readdata;
  wire             std_2s60_burst_8_downstream_readdatavalid;
  wire             std_2s60_burst_8_downstream_reset_n;
  wire             std_2s60_burst_8_downstream_run;
  wire             std_2s60_burst_8_downstream_waitrequest;
  reg              std_2s60_burst_8_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_8_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_8_downstream_requests_lan91c111_s1) & (std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_8_downstream_requests_ext_ram_s1) & (std_2s60_burst_8_downstream_granted_lan91c111_s1 | ~std_2s60_burst_8_downstream_qualified_request_lan91c111_s1) & (std_2s60_burst_8_downstream_granted_ext_ram_s1 | ~std_2s60_burst_8_downstream_qualified_request_ext_ram_s1) & ((~std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_8_downstream_read | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_8_downstream_read))) & ((~std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_8_downstream_write | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_8_downstream_write))) & ((~std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_8_downstream_read | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_8_downstream_read))) & ((~std_2s60_burst_8_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_8_downstream_write | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_8_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_8_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_8_downstream_address_to_slave = std_2s60_burst_8_downstream_address;

  //std_2s60_burst_8_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_8_downstream_read_but_no_slave_selected <= std_2s60_burst_8_downstream_read & std_2s60_burst_8_downstream_run & ~std_2s60_burst_8_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_8_downstream_is_granted_some_slave = std_2s60_burst_8_downstream_granted_lan91c111_s1 |
    std_2s60_burst_8_downstream_granted_ext_ram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_8_downstream_readdatavalid = std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1 |
    std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_8_downstream_readdatavalid = std_2s60_burst_8_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_8_downstream_readdatavalid |
    std_2s60_burst_8_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_8_downstream_readdatavalid;

  //std_2s60_burst_8/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_8_downstream_readdata = ({32 {~std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1}} | incoming_ext_ram_bus_data) &
    ({32 {~std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1}} | incoming_ext_ram_bus_data);

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_8_downstream_waitrequest = ~std_2s60_burst_8_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_8_downstream_latency_counter <= p1_std_2s60_burst_8_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_8_downstream_latency_counter = ((std_2s60_burst_8_downstream_run & std_2s60_burst_8_downstream_read))? latency_load_value :
    (std_2s60_burst_8_downstream_latency_counter)? std_2s60_burst_8_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {std_2s60_burst_8_downstream_requests_lan91c111_s1}} & 2) |
    ({2 {std_2s60_burst_8_downstream_requests_ext_ram_s1}} & 2);

  //std_2s60_burst_8_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_8_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_8_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_address_last_time <= std_2s60_burst_8_downstream_address;
    end


  //std_2s60_burst_8/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_8_downstream_waitrequest & (std_2s60_burst_8_downstream_read | std_2s60_burst_8_downstream_write);
    end


  //std_2s60_burst_8_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_address != std_2s60_burst_8_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_8_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_burstcount_last_time <= std_2s60_burst_8_downstream_burstcount;
    end


  //std_2s60_burst_8_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_burstcount != std_2s60_burst_8_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_8_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_byteenable_last_time <= std_2s60_burst_8_downstream_byteenable;
    end


  //std_2s60_burst_8_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_byteenable != std_2s60_burst_8_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_8_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_read_last_time <= std_2s60_burst_8_downstream_read;
    end


  //std_2s60_burst_8_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_read != std_2s60_burst_8_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_8_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_write_last_time <= std_2s60_burst_8_downstream_write;
    end


  //std_2s60_burst_8_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_write != std_2s60_burst_8_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_8_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_8_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_8_downstream_writedata_last_time <= std_2s60_burst_8_downstream_writedata;
    end


  //std_2s60_burst_8_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_8_downstream_writedata != std_2s60_burst_8_downstream_writedata_last_time) & std_2s60_burst_8_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_8_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_std_2s60_burst_9_upstream_module (
                                                              // inputs:
                                                               clear_fifo,
                                                               clk,
                                                               data_in,
                                                               read,
                                                               reset_n,
                                                               sync_reset,
                                                               write,

                                                              // outputs:
                                                               data_out,
                                                               empty,
                                                               fifo_contains_ones_n,
                                                               full
                                                            )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_9_upstream_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_9_upstream_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_burstcount,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_debugaccess,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register,
                                               cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register,
                                               cpu_data_master_write,
                                               cpu_data_master_writedata,
                                               reset_n,
                                               std_2s60_burst_9_upstream_readdata,
                                               std_2s60_burst_9_upstream_readdatavalid,
                                               std_2s60_burst_9_upstream_waitrequest,

                                              // outputs:
                                               cpu_data_master_granted_std_2s60_burst_9_upstream,
                                               cpu_data_master_qualified_request_std_2s60_burst_9_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream,
                                               cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register,
                                               cpu_data_master_requests_std_2s60_burst_9_upstream,
                                               d1_std_2s60_burst_9_upstream_end_xfer,
                                               std_2s60_burst_9_upstream_address,
                                               std_2s60_burst_9_upstream_burstcount,
                                               std_2s60_burst_9_upstream_byteaddress,
                                               std_2s60_burst_9_upstream_byteenable,
                                               std_2s60_burst_9_upstream_debugaccess,
                                               std_2s60_burst_9_upstream_read,
                                               std_2s60_burst_9_upstream_readdata_from_sa,
                                               std_2s60_burst_9_upstream_waitrequest_from_sa,
                                               std_2s60_burst_9_upstream_write,
                                               std_2s60_burst_9_upstream_writedata
                                            )
;

  output           cpu_data_master_granted_std_2s60_burst_9_upstream;
  output           cpu_data_master_qualified_request_std_2s60_burst_9_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_9_upstream;
  output           cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  output           cpu_data_master_requests_std_2s60_burst_9_upstream;
  output           d1_std_2s60_burst_9_upstream_end_xfer;
  output  [ 15: 0] std_2s60_burst_9_upstream_address;
  output  [  3: 0] std_2s60_burst_9_upstream_burstcount;
  output  [ 17: 0] std_2s60_burst_9_upstream_byteaddress;
  output  [  3: 0] std_2s60_burst_9_upstream_byteenable;
  output           std_2s60_burst_9_upstream_debugaccess;
  output           std_2s60_burst_9_upstream_read;
  output  [ 31: 0] std_2s60_burst_9_upstream_readdata_from_sa;
  output           std_2s60_burst_9_upstream_waitrequest_from_sa;
  output           std_2s60_burst_9_upstream_write;
  output  [ 31: 0] std_2s60_burst_9_upstream_writedata;
  input            clk;
  input   [ 25: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  input            cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] std_2s60_burst_9_upstream_readdata;
  input            std_2s60_burst_9_upstream_readdatavalid;
  input            std_2s60_burst_9_upstream_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_std_2s60_burst_9_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_9_upstream;
  wire             cpu_data_master_rdv_fifo_empty_std_2s60_burst_9_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_std_2s60_burst_9_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_9_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  wire             cpu_data_master_requests_std_2s60_burst_9_upstream;
  wire             cpu_data_master_saved_grant_std_2s60_burst_9_upstream;
  reg              d1_reasons_to_wait;
  reg              d1_std_2s60_burst_9_upstream_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_std_2s60_burst_9_upstream_load_fifo;
  wire    [ 25: 0] shifted_address_to_std_2s60_burst_9_upstream_from_cpu_data_master;
  wire    [ 15: 0] std_2s60_burst_9_upstream_address;
  wire             std_2s60_burst_9_upstream_allgrants;
  wire             std_2s60_burst_9_upstream_allow_new_arb_cycle;
  wire             std_2s60_burst_9_upstream_any_bursting_master_saved_grant;
  wire             std_2s60_burst_9_upstream_any_continuerequest;
  wire             std_2s60_burst_9_upstream_arb_counter_enable;
  reg     [  7: 0] std_2s60_burst_9_upstream_arb_share_counter;
  wire    [  7: 0] std_2s60_burst_9_upstream_arb_share_counter_next_value;
  wire    [  7: 0] std_2s60_burst_9_upstream_arb_share_set_values;
  reg     [  2: 0] std_2s60_burst_9_upstream_bbt_burstcounter;
  wire             std_2s60_burst_9_upstream_beginbursttransfer_internal;
  wire             std_2s60_burst_9_upstream_begins_xfer;
  wire    [  3: 0] std_2s60_burst_9_upstream_burstcount;
  wire             std_2s60_burst_9_upstream_burstcount_fifo_empty;
  wire    [ 17: 0] std_2s60_burst_9_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_9_upstream_byteenable;
  reg     [  3: 0] std_2s60_burst_9_upstream_current_burst;
  wire    [  3: 0] std_2s60_burst_9_upstream_current_burst_minus_one;
  wire             std_2s60_burst_9_upstream_debugaccess;
  wire             std_2s60_burst_9_upstream_end_xfer;
  wire             std_2s60_burst_9_upstream_firsttransfer;
  wire             std_2s60_burst_9_upstream_grant_vector;
  wire             std_2s60_burst_9_upstream_in_a_read_cycle;
  wire             std_2s60_burst_9_upstream_in_a_write_cycle;
  reg              std_2s60_burst_9_upstream_load_fifo;
  wire             std_2s60_burst_9_upstream_master_qreq_vector;
  wire             std_2s60_burst_9_upstream_move_on_to_next_transaction;
  wire    [  2: 0] std_2s60_burst_9_upstream_next_bbt_burstcount;
  wire    [  3: 0] std_2s60_burst_9_upstream_next_burst_count;
  wire             std_2s60_burst_9_upstream_non_bursting_master_requests;
  wire             std_2s60_burst_9_upstream_read;
  wire    [ 31: 0] std_2s60_burst_9_upstream_readdata_from_sa;
  wire             std_2s60_burst_9_upstream_readdatavalid_from_sa;
  reg              std_2s60_burst_9_upstream_reg_firsttransfer;
  wire    [  3: 0] std_2s60_burst_9_upstream_selected_burstcount;
  reg              std_2s60_burst_9_upstream_slavearbiterlockenable;
  wire             std_2s60_burst_9_upstream_slavearbiterlockenable2;
  wire             std_2s60_burst_9_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] std_2s60_burst_9_upstream_transaction_burst_count;
  wire             std_2s60_burst_9_upstream_unreg_firsttransfer;
  wire             std_2s60_burst_9_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_9_upstream_waits_for_read;
  wire             std_2s60_burst_9_upstream_waits_for_write;
  wire             std_2s60_burst_9_upstream_write;
  wire    [ 31: 0] std_2s60_burst_9_upstream_writedata;
  wire             wait_for_std_2s60_burst_9_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~std_2s60_burst_9_upstream_end_xfer;
    end


  assign std_2s60_burst_9_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_std_2s60_burst_9_upstream));
  //assign std_2s60_burst_9_upstream_readdatavalid_from_sa = std_2s60_burst_9_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_9_upstream_readdatavalid_from_sa = std_2s60_burst_9_upstream_readdatavalid;

  //assign std_2s60_burst_9_upstream_readdata_from_sa = std_2s60_burst_9_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_9_upstream_readdata_from_sa = std_2s60_burst_9_upstream_readdata;

  assign cpu_data_master_requests_std_2s60_burst_9_upstream = ({cpu_data_master_address_to_slave[25 : 16] , 16'b0} == 26'h2110000) & (cpu_data_master_read | cpu_data_master_write);
  //assign std_2s60_burst_9_upstream_waitrequest_from_sa = std_2s60_burst_9_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign std_2s60_burst_9_upstream_waitrequest_from_sa = std_2s60_burst_9_upstream_waitrequest;

  //std_2s60_burst_9_upstream_arb_share_counter set values, which is an e_mux
  assign std_2s60_burst_9_upstream_arb_share_set_values = (cpu_data_master_granted_std_2s60_burst_9_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //std_2s60_burst_9_upstream_non_bursting_master_requests mux, which is an e_mux
  assign std_2s60_burst_9_upstream_non_bursting_master_requests = 0;

  //std_2s60_burst_9_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign std_2s60_burst_9_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_std_2s60_burst_9_upstream;

  //std_2s60_burst_9_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign std_2s60_burst_9_upstream_arb_share_counter_next_value = std_2s60_burst_9_upstream_firsttransfer ? (std_2s60_burst_9_upstream_arb_share_set_values - 1) : |std_2s60_burst_9_upstream_arb_share_counter ? (std_2s60_burst_9_upstream_arb_share_counter - 1) : 0;

  //std_2s60_burst_9_upstream_allgrants all slave grants, which is an e_mux
  assign std_2s60_burst_9_upstream_allgrants = |std_2s60_burst_9_upstream_grant_vector;

  //std_2s60_burst_9_upstream_end_xfer assignment, which is an e_assign
  assign std_2s60_burst_9_upstream_end_xfer = ~(std_2s60_burst_9_upstream_waits_for_read | std_2s60_burst_9_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream = std_2s60_burst_9_upstream_end_xfer & (~std_2s60_burst_9_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //std_2s60_burst_9_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign std_2s60_burst_9_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream & std_2s60_burst_9_upstream_allgrants) | (end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream & ~std_2s60_burst_9_upstream_non_bursting_master_requests);

  //std_2s60_burst_9_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_arb_share_counter <= 0;
      else if (std_2s60_burst_9_upstream_arb_counter_enable)
          std_2s60_burst_9_upstream_arb_share_counter <= std_2s60_burst_9_upstream_arb_share_counter_next_value;
    end


  //std_2s60_burst_9_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_slavearbiterlockenable <= 0;
      else if ((|std_2s60_burst_9_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream) | (end_xfer_arb_share_counter_term_std_2s60_burst_9_upstream & ~std_2s60_burst_9_upstream_non_bursting_master_requests))
          std_2s60_burst_9_upstream_slavearbiterlockenable <= |std_2s60_burst_9_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master std_2s60_burst_9/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = std_2s60_burst_9_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //std_2s60_burst_9_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign std_2s60_burst_9_upstream_slavearbiterlockenable2 = |std_2s60_burst_9_upstream_arb_share_counter_next_value;

  //cpu/data_master std_2s60_burst_9/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = std_2s60_burst_9_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //std_2s60_burst_9_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign std_2s60_burst_9_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_std_2s60_burst_9_upstream = cpu_data_master_requests_std_2s60_burst_9_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register) | (|cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register))));
  //unique name for std_2s60_burst_9_upstream_move_on_to_next_transaction, which is an e_assign
  assign std_2s60_burst_9_upstream_move_on_to_next_transaction = std_2s60_burst_9_upstream_this_cycle_is_the_last_burst & std_2s60_burst_9_upstream_load_fifo;

  //the currently selected burstcount for std_2s60_burst_9_upstream, which is an e_mux
  assign std_2s60_burst_9_upstream_selected_burstcount = (cpu_data_master_granted_std_2s60_burst_9_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_std_2s60_burst_9_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_std_2s60_burst_9_upstream_module burstcount_fifo_for_std_2s60_burst_9_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (std_2s60_burst_9_upstream_selected_burstcount),
      .data_out             (std_2s60_burst_9_upstream_transaction_burst_count),
      .empty                (std_2s60_burst_9_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (std_2s60_burst_9_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read & std_2s60_burst_9_upstream_load_fifo & ~(std_2s60_burst_9_upstream_this_cycle_is_the_last_burst & std_2s60_burst_9_upstream_burstcount_fifo_empty))
    );

  //std_2s60_burst_9_upstream current burst minus one, which is an e_assign
  assign std_2s60_burst_9_upstream_current_burst_minus_one = std_2s60_burst_9_upstream_current_burst - 1;

  //what to load in current_burst, for std_2s60_burst_9_upstream, which is an e_mux
  assign std_2s60_burst_9_upstream_next_burst_count = (((in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read) & ~std_2s60_burst_9_upstream_load_fifo))? std_2s60_burst_9_upstream_selected_burstcount :
    ((in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read & std_2s60_burst_9_upstream_this_cycle_is_the_last_burst & std_2s60_burst_9_upstream_burstcount_fifo_empty))? std_2s60_burst_9_upstream_selected_burstcount :
    (std_2s60_burst_9_upstream_this_cycle_is_the_last_burst)? std_2s60_burst_9_upstream_transaction_burst_count :
    std_2s60_burst_9_upstream_current_burst_minus_one;

  //the current burst count for std_2s60_burst_9_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_current_burst <= 0;
      else if (std_2s60_burst_9_upstream_readdatavalid_from_sa | (~std_2s60_burst_9_upstream_load_fifo & (in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read)))
          std_2s60_burst_9_upstream_current_burst <= std_2s60_burst_9_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_std_2s60_burst_9_upstream_load_fifo = (~std_2s60_burst_9_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read) & std_2s60_burst_9_upstream_load_fifo))? 1 :
    ~std_2s60_burst_9_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read) & ~std_2s60_burst_9_upstream_load_fifo | std_2s60_burst_9_upstream_this_cycle_is_the_last_burst)
          std_2s60_burst_9_upstream_load_fifo <= p0_std_2s60_burst_9_upstream_load_fifo;
    end


  //the last cycle in the burst for std_2s60_burst_9_upstream, which is an e_assign
  assign std_2s60_burst_9_upstream_this_cycle_is_the_last_burst = ~(|std_2s60_burst_9_upstream_current_burst_minus_one) & std_2s60_burst_9_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_std_2s60_burst_9_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_std_2s60_burst_9_upstream_module rdv_fifo_for_cpu_data_master_to_std_2s60_burst_9_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_std_2s60_burst_9_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_std_2s60_burst_9_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_std_2s60_burst_9_upstream),
      .full                 (),
      .read                 (std_2s60_burst_9_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~std_2s60_burst_9_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_std_2s60_burst_9_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_std_2s60_burst_9_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_std_2s60_burst_9_upstream = std_2s60_burst_9_upstream_readdatavalid_from_sa;

  //std_2s60_burst_9_upstream_writedata mux, which is an e_mux
  assign std_2s60_burst_9_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for std_2s60_burst_9/upstream, which is an e_mux
  assign std_2s60_burst_9_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_std_2s60_burst_9_upstream = cpu_data_master_qualified_request_std_2s60_burst_9_upstream;

  //cpu/data_master saved-grant std_2s60_burst_9/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_std_2s60_burst_9_upstream = cpu_data_master_requests_std_2s60_burst_9_upstream;

  //allow new arb cycle for std_2s60_burst_9/upstream, which is an e_assign
  assign std_2s60_burst_9_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign std_2s60_burst_9_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign std_2s60_burst_9_upstream_master_qreq_vector = 1;

  //std_2s60_burst_9_upstream_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_9_upstream_firsttransfer = std_2s60_burst_9_upstream_begins_xfer ? std_2s60_burst_9_upstream_unreg_firsttransfer : std_2s60_burst_9_upstream_reg_firsttransfer;

  //std_2s60_burst_9_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign std_2s60_burst_9_upstream_unreg_firsttransfer = ~(std_2s60_burst_9_upstream_slavearbiterlockenable & std_2s60_burst_9_upstream_any_continuerequest);

  //std_2s60_burst_9_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_reg_firsttransfer <= 1'b1;
      else if (std_2s60_burst_9_upstream_begins_xfer)
          std_2s60_burst_9_upstream_reg_firsttransfer <= std_2s60_burst_9_upstream_unreg_firsttransfer;
    end


  //std_2s60_burst_9_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign std_2s60_burst_9_upstream_next_bbt_burstcount = ((((std_2s60_burst_9_upstream_write) && (std_2s60_burst_9_upstream_bbt_burstcounter == 0))))? (std_2s60_burst_9_upstream_burstcount - 1) :
    ((((std_2s60_burst_9_upstream_read) && (std_2s60_burst_9_upstream_bbt_burstcounter == 0))))? 0 :
    (std_2s60_burst_9_upstream_bbt_burstcounter - 1);

  //std_2s60_burst_9_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_upstream_bbt_burstcounter <= 0;
      else if (std_2s60_burst_9_upstream_begins_xfer)
          std_2s60_burst_9_upstream_bbt_burstcounter <= std_2s60_burst_9_upstream_next_bbt_burstcount;
    end


  //std_2s60_burst_9_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign std_2s60_burst_9_upstream_beginbursttransfer_internal = std_2s60_burst_9_upstream_begins_xfer & (std_2s60_burst_9_upstream_bbt_burstcounter == 0);

  //std_2s60_burst_9_upstream_read assignment, which is an e_mux
  assign std_2s60_burst_9_upstream_read = cpu_data_master_granted_std_2s60_burst_9_upstream & cpu_data_master_read;

  //std_2s60_burst_9_upstream_write assignment, which is an e_mux
  assign std_2s60_burst_9_upstream_write = cpu_data_master_granted_std_2s60_burst_9_upstream & cpu_data_master_write;

  assign shifted_address_to_std_2s60_burst_9_upstream_from_cpu_data_master = cpu_data_master_address_to_slave;
  //std_2s60_burst_9_upstream_address mux, which is an e_mux
  assign std_2s60_burst_9_upstream_address = shifted_address_to_std_2s60_burst_9_upstream_from_cpu_data_master >> 2;

  //d1_std_2s60_burst_9_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_std_2s60_burst_9_upstream_end_xfer <= 1;
      else if (1)
          d1_std_2s60_burst_9_upstream_end_xfer <= std_2s60_burst_9_upstream_end_xfer;
    end


  //std_2s60_burst_9_upstream_waits_for_read in a cycle, which is an e_mux
  assign std_2s60_burst_9_upstream_waits_for_read = std_2s60_burst_9_upstream_in_a_read_cycle & std_2s60_burst_9_upstream_waitrequest_from_sa;

  //std_2s60_burst_9_upstream_in_a_read_cycle assignment, which is an e_assign
  assign std_2s60_burst_9_upstream_in_a_read_cycle = cpu_data_master_granted_std_2s60_burst_9_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = std_2s60_burst_9_upstream_in_a_read_cycle;

  //std_2s60_burst_9_upstream_waits_for_write in a cycle, which is an e_mux
  assign std_2s60_burst_9_upstream_waits_for_write = std_2s60_burst_9_upstream_in_a_write_cycle & std_2s60_burst_9_upstream_waitrequest_from_sa;

  //std_2s60_burst_9_upstream_in_a_write_cycle assignment, which is an e_assign
  assign std_2s60_burst_9_upstream_in_a_write_cycle = cpu_data_master_granted_std_2s60_burst_9_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = std_2s60_burst_9_upstream_in_a_write_cycle;

  assign wait_for_std_2s60_burst_9_upstream_counter = 0;
  //std_2s60_burst_9_upstream_byteenable byte enable port mux, which is an e_mux
  assign std_2s60_burst_9_upstream_byteenable = (cpu_data_master_granted_std_2s60_burst_9_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign std_2s60_burst_9_upstream_burstcount = (cpu_data_master_granted_std_2s60_burst_9_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign std_2s60_burst_9_upstream_debugaccess = (cpu_data_master_granted_std_2s60_burst_9_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_9/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_std_2s60_burst_9_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave std_2s60_burst_9/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_burst_9_downstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 d1_ext_ram_bus_avalon_slave_end_xfer,
                                                 ext_ram_s1_wait_counter_eq_0,
                                                 incoming_ext_ram_bus_data,
                                                 lan91c111_s1_wait_counter_eq_0,
                                                 reset_n,
                                                 std_2s60_burst_9_downstream_address,
                                                 std_2s60_burst_9_downstream_burstcount,
                                                 std_2s60_burst_9_downstream_byteenable,
                                                 std_2s60_burst_9_downstream_granted_ext_ram_s1,
                                                 std_2s60_burst_9_downstream_granted_lan91c111_s1,
                                                 std_2s60_burst_9_downstream_qualified_request_ext_ram_s1,
                                                 std_2s60_burst_9_downstream_qualified_request_lan91c111_s1,
                                                 std_2s60_burst_9_downstream_read,
                                                 std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1,
                                                 std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1,
                                                 std_2s60_burst_9_downstream_requests_ext_ram_s1,
                                                 std_2s60_burst_9_downstream_requests_lan91c111_s1,
                                                 std_2s60_burst_9_downstream_write,
                                                 std_2s60_burst_9_downstream_writedata,

                                                // outputs:
                                                 std_2s60_burst_9_downstream_address_to_slave,
                                                 std_2s60_burst_9_downstream_latency_counter,
                                                 std_2s60_burst_9_downstream_readdata,
                                                 std_2s60_burst_9_downstream_readdatavalid,
                                                 std_2s60_burst_9_downstream_reset_n,
                                                 std_2s60_burst_9_downstream_waitrequest
                                              )
;

  output  [ 15: 0] std_2s60_burst_9_downstream_address_to_slave;
  output  [  1: 0] std_2s60_burst_9_downstream_latency_counter;
  output  [ 31: 0] std_2s60_burst_9_downstream_readdata;
  output           std_2s60_burst_9_downstream_readdatavalid;
  output           std_2s60_burst_9_downstream_reset_n;
  output           std_2s60_burst_9_downstream_waitrequest;
  input            clk;
  input            d1_ext_ram_bus_avalon_slave_end_xfer;
  input            ext_ram_s1_wait_counter_eq_0;
  input   [ 31: 0] incoming_ext_ram_bus_data;
  input            lan91c111_s1_wait_counter_eq_0;
  input            reset_n;
  input   [ 15: 0] std_2s60_burst_9_downstream_address;
  input            std_2s60_burst_9_downstream_burstcount;
  input   [  3: 0] std_2s60_burst_9_downstream_byteenable;
  input            std_2s60_burst_9_downstream_granted_ext_ram_s1;
  input            std_2s60_burst_9_downstream_granted_lan91c111_s1;
  input            std_2s60_burst_9_downstream_qualified_request_ext_ram_s1;
  input            std_2s60_burst_9_downstream_qualified_request_lan91c111_s1;
  input            std_2s60_burst_9_downstream_read;
  input            std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1;
  input            std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1;
  input            std_2s60_burst_9_downstream_requests_ext_ram_s1;
  input            std_2s60_burst_9_downstream_requests_lan91c111_s1;
  input            std_2s60_burst_9_downstream_write;
  input   [ 31: 0] std_2s60_burst_9_downstream_writedata;

  reg              active_and_waiting_last_time;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] p1_std_2s60_burst_9_downstream_latency_counter;
  wire             pre_flush_std_2s60_burst_9_downstream_readdatavalid;
  wire             r_0;
  reg     [ 15: 0] std_2s60_burst_9_downstream_address_last_time;
  wire    [ 15: 0] std_2s60_burst_9_downstream_address_to_slave;
  reg              std_2s60_burst_9_downstream_burstcount_last_time;
  reg     [  3: 0] std_2s60_burst_9_downstream_byteenable_last_time;
  wire             std_2s60_burst_9_downstream_is_granted_some_slave;
  reg     [  1: 0] std_2s60_burst_9_downstream_latency_counter;
  reg              std_2s60_burst_9_downstream_read_but_no_slave_selected;
  reg              std_2s60_burst_9_downstream_read_last_time;
  wire    [ 31: 0] std_2s60_burst_9_downstream_readdata;
  wire             std_2s60_burst_9_downstream_readdatavalid;
  wire             std_2s60_burst_9_downstream_reset_n;
  wire             std_2s60_burst_9_downstream_run;
  wire             std_2s60_burst_9_downstream_waitrequest;
  reg              std_2s60_burst_9_downstream_write_last_time;
  reg     [ 31: 0] std_2s60_burst_9_downstream_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_9_downstream_requests_lan91c111_s1) & (std_2s60_burst_9_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_9_downstream_requests_ext_ram_s1) & (std_2s60_burst_9_downstream_granted_lan91c111_s1 | ~std_2s60_burst_9_downstream_qualified_request_lan91c111_s1) & (std_2s60_burst_9_downstream_granted_ext_ram_s1 | ~std_2s60_burst_9_downstream_qualified_request_ext_ram_s1) & ((~std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_9_downstream_read | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_9_downstream_read))) & ((~std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 | ~std_2s60_burst_9_downstream_write | (1 & ((lan91c111_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_9_downstream_write))) & ((~std_2s60_burst_9_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_9_downstream_read | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_9_downstream_read))) & ((~std_2s60_burst_9_downstream_qualified_request_ext_ram_s1 | ~std_2s60_burst_9_downstream_write | (1 & ((ext_ram_s1_wait_counter_eq_0 & ~d1_ext_ram_bus_avalon_slave_end_xfer)) & std_2s60_burst_9_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign std_2s60_burst_9_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign std_2s60_burst_9_downstream_address_to_slave = std_2s60_burst_9_downstream_address;

  //std_2s60_burst_9_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_read_but_no_slave_selected <= 0;
      else if (1)
          std_2s60_burst_9_downstream_read_but_no_slave_selected <= std_2s60_burst_9_downstream_read & std_2s60_burst_9_downstream_run & ~std_2s60_burst_9_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign std_2s60_burst_9_downstream_is_granted_some_slave = std_2s60_burst_9_downstream_granted_lan91c111_s1 |
    std_2s60_burst_9_downstream_granted_ext_ram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_std_2s60_burst_9_downstream_readdatavalid = std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1 |
    std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign std_2s60_burst_9_downstream_readdatavalid = std_2s60_burst_9_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_9_downstream_readdatavalid |
    std_2s60_burst_9_downstream_read_but_no_slave_selected |
    pre_flush_std_2s60_burst_9_downstream_readdatavalid;

  //std_2s60_burst_9/downstream readdata mux, which is an e_mux
  assign std_2s60_burst_9_downstream_readdata = ({32 {~std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1}} | incoming_ext_ram_bus_data) &
    ({32 {~std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1}} | incoming_ext_ram_bus_data);

  //actual waitrequest port, which is an e_assign
  assign std_2s60_burst_9_downstream_waitrequest = ~std_2s60_burst_9_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_latency_counter <= 0;
      else if (1)
          std_2s60_burst_9_downstream_latency_counter <= p1_std_2s60_burst_9_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_std_2s60_burst_9_downstream_latency_counter = ((std_2s60_burst_9_downstream_run & std_2s60_burst_9_downstream_read))? latency_load_value :
    (std_2s60_burst_9_downstream_latency_counter)? std_2s60_burst_9_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {std_2s60_burst_9_downstream_requests_lan91c111_s1}} & 2) |
    ({2 {std_2s60_burst_9_downstream_requests_ext_ram_s1}} & 2);

  //std_2s60_burst_9_downstream_reset_n assignment, which is an e_assign
  assign std_2s60_burst_9_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //std_2s60_burst_9_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_address_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_address_last_time <= std_2s60_burst_9_downstream_address;
    end


  //std_2s60_burst_9/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else if (1)
          active_and_waiting_last_time <= std_2s60_burst_9_downstream_waitrequest & (std_2s60_burst_9_downstream_read | std_2s60_burst_9_downstream_write);
    end


  //std_2s60_burst_9_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_address != std_2s60_burst_9_downstream_address_last_time))
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_9_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_burstcount_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_burstcount_last_time <= std_2s60_burst_9_downstream_burstcount;
    end


  //std_2s60_burst_9_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_burstcount != std_2s60_burst_9_downstream_burstcount_last_time))
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_9_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_byteenable_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_byteenable_last_time <= std_2s60_burst_9_downstream_byteenable;
    end


  //std_2s60_burst_9_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_byteenable != std_2s60_burst_9_downstream_byteenable_last_time))
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_9_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_read_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_read_last_time <= std_2s60_burst_9_downstream_read;
    end


  //std_2s60_burst_9_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_read != std_2s60_burst_9_downstream_read_last_time))
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_9_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_write_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_write_last_time <= std_2s60_burst_9_downstream_write;
    end


  //std_2s60_burst_9_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_write != std_2s60_burst_9_downstream_write_last_time))
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //std_2s60_burst_9_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          std_2s60_burst_9_downstream_writedata_last_time <= 0;
      else if (1)
          std_2s60_burst_9_downstream_writedata_last_time <= std_2s60_burst_9_downstream_writedata;
    end


  //std_2s60_burst_9_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (std_2s60_burst_9_downstream_writedata != std_2s60_burst_9_downstream_writedata_last_time) & std_2s60_burst_9_downstream_write)
        begin
          $write("%0d ns: std_2s60_burst_9_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sys_clk_timer_s1_arbitrator (
                                     // inputs:
                                      clk,
                                      reset_n,
                                      std_2s60_burst_10_downstream_address_to_slave,
                                      std_2s60_burst_10_downstream_arbitrationshare,
                                      std_2s60_burst_10_downstream_burstcount,
                                      std_2s60_burst_10_downstream_latency_counter,
                                      std_2s60_burst_10_downstream_nativeaddress,
                                      std_2s60_burst_10_downstream_read,
                                      std_2s60_burst_10_downstream_write,
                                      std_2s60_burst_10_downstream_writedata,
                                      sys_clk_timer_s1_irq,
                                      sys_clk_timer_s1_readdata,

                                     // outputs:
                                      d1_sys_clk_timer_s1_end_xfer,
                                      std_2s60_burst_10_downstream_granted_sys_clk_timer_s1,
                                      std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1,
                                      std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1,
                                      std_2s60_burst_10_downstream_requests_sys_clk_timer_s1,
                                      sys_clk_timer_s1_address,
                                      sys_clk_timer_s1_chipselect,
                                      sys_clk_timer_s1_irq_from_sa,
                                      sys_clk_timer_s1_readdata_from_sa,
                                      sys_clk_timer_s1_reset_n,
                                      sys_clk_timer_s1_write_n,
                                      sys_clk_timer_s1_writedata
                                   )
;

  output           d1_sys_clk_timer_s1_end_xfer;
  output           std_2s60_burst_10_downstream_granted_sys_clk_timer_s1;
  output           std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1;
  output           std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1;
  output           std_2s60_burst_10_downstream_requests_sys_clk_timer_s1;
  output  [  2: 0] sys_clk_timer_s1_address;
  output           sys_clk_timer_s1_chipselect;
  output           sys_clk_timer_s1_irq_from_sa;
  output  [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  output           sys_clk_timer_s1_reset_n;
  output           sys_clk_timer_s1_write_n;
  output  [ 15: 0] sys_clk_timer_s1_writedata;
  input            clk;
  input            reset_n;
  input   [  3: 0] std_2s60_burst_10_downstream_address_to_slave;
  input   [  4: 0] std_2s60_burst_10_downstream_arbitrationshare;
  input            std_2s60_burst_10_downstream_burstcount;
  input            std_2s60_burst_10_downstream_latency_counter;
  input   [  3: 0] std_2s60_burst_10_downstream_nativeaddress;
  input            std_2s60_burst_10_downstream_read;
  input            std_2s60_burst_10_downstream_write;
  input   [ 15: 0] std_2s60_burst_10_downstream_writedata;
  input            sys_clk_timer_s1_irq;
  input   [ 15: 0] sys_clk_timer_s1_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sys_clk_timer_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sys_clk_timer_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             std_2s60_burst_10_downstream_arbiterlock;
  wire             std_2s60_burst_10_downstream_arbiterlock2;
  wire             std_2s60_burst_10_downstream_continuerequest;
  wire             std_2s60_burst_10_downstream_granted_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_requests_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_saved_grant_sys_clk_timer_s1;
  wire    [  2: 0] sys_clk_timer_s1_address;
  wire             sys_clk_timer_s1_allgrants;
  wire             sys_clk_timer_s1_allow_new_arb_cycle;
  wire             sys_clk_timer_s1_any_bursting_master_saved_grant;
  wire             sys_clk_timer_s1_any_continuerequest;
  wire             sys_clk_timer_s1_arb_counter_enable;
  reg     [  4: 0] sys_clk_timer_s1_arb_share_counter;
  wire    [  4: 0] sys_clk_timer_s1_arb_share_counter_next_value;
  wire    [  4: 0] sys_clk_timer_s1_arb_share_set_values;
  wire             sys_clk_timer_s1_beginbursttransfer_internal;
  wire             sys_clk_timer_s1_begins_xfer;
  wire             sys_clk_timer_s1_chipselect;
  wire             sys_clk_timer_s1_end_xfer;
  wire             sys_clk_timer_s1_firsttransfer;
  wire             sys_clk_timer_s1_grant_vector;
  wire             sys_clk_timer_s1_in_a_read_cycle;
  wire             sys_clk_timer_s1_in_a_write_cycle;
  wire             sys_clk_timer_s1_irq_from_sa;
  wire             sys_clk_timer_s1_master_qreq_vector;
  wire             sys_clk_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  reg              sys_clk_timer_s1_reg_firsttransfer;
  wire             sys_clk_timer_s1_reset_n;
  reg              sys_clk_timer_s1_slavearbiterlockenable;
  wire             sys_clk_timer_s1_slavearbiterlockenable2;
  wire             sys_clk_timer_s1_unreg_firsttransfer;
  wire             sys_clk_timer_s1_waits_for_read;
  wire             sys_clk_timer_s1_waits_for_write;
  wire             sys_clk_timer_s1_write_n;
  wire    [ 15: 0] sys_clk_timer_s1_writedata;
  wire             wait_for_sys_clk_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~sys_clk_timer_s1_end_xfer;
    end


  assign sys_clk_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1));
  //assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata;

  assign std_2s60_burst_10_downstream_requests_sys_clk_timer_s1 = (1) & (std_2s60_burst_10_downstream_read | std_2s60_burst_10_downstream_write);
  //sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  assign sys_clk_timer_s1_arb_share_set_values = (std_2s60_burst_10_downstream_granted_sys_clk_timer_s1)? std_2s60_burst_10_downstream_arbitrationshare :
    1;

  //sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign sys_clk_timer_s1_non_bursting_master_requests = 0;

  //sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sys_clk_timer_s1_any_bursting_master_saved_grant = std_2s60_burst_10_downstream_saved_grant_sys_clk_timer_s1;

  //sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sys_clk_timer_s1_arb_share_counter_next_value = sys_clk_timer_s1_firsttransfer ? (sys_clk_timer_s1_arb_share_set_values - 1) : |sys_clk_timer_s1_arb_share_counter ? (sys_clk_timer_s1_arb_share_counter - 1) : 0;

  //sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  assign sys_clk_timer_s1_allgrants = |sys_clk_timer_s1_grant_vector;

  //sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  assign sys_clk_timer_s1_end_xfer = ~(sys_clk_timer_s1_waits_for_read | sys_clk_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sys_clk_timer_s1 = sys_clk_timer_s1_end_xfer & (~sys_clk_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sys_clk_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & sys_clk_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & ~sys_clk_timer_s1_non_bursting_master_requests);

  //sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_arb_share_counter <= 0;
      else if (sys_clk_timer_s1_arb_counter_enable)
          sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
    end


  //sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_slavearbiterlockenable <= 0;
      else if ((|sys_clk_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sys_clk_timer_s1) | (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & ~sys_clk_timer_s1_non_bursting_master_requests))
          sys_clk_timer_s1_slavearbiterlockenable <= |sys_clk_timer_s1_arb_share_counter_next_value;
    end


  //std_2s60_burst_10/downstream sys_clk_timer/s1 arbiterlock, which is an e_assign
  assign std_2s60_burst_10_downstream_arbiterlock = sys_clk_timer_s1_slavearbiterlockenable & std_2s60_burst_10_downstream_continuerequest;

  //sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sys_clk_timer_s1_slavearbiterlockenable2 = |sys_clk_timer_s1_arb_share_counter_next_value;

  //std_2s60_burst_10/downstream sys_clk_timer/s1 arbiterlock2, which is an e_assign
  assign std_2s60_burst_10_downstream_arbiterlock2 = sys_clk_timer_s1_slavearbiterlockenable2 & std_2s60_burst_10_downstream_continuerequest;

  //sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sys_clk_timer_s1_any_continuerequest = 1;

  //std_2s60_burst_10_downstream_continuerequest continued request, which is an e_assign
  assign std_2s60_burst_10_downstream_continuerequest = 1;

  assign std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 = std_2s60_burst_10_downstream_requests_sys_clk_timer_s1 & ~((std_2s60_burst_10_downstream_read & ((std_2s60_burst_10_downstream_latency_counter != 0))));
  //local readdatavalid std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1, which is an e_mux
  assign std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1 = std_2s60_burst_10_downstream_granted_sys_clk_timer_s1 & std_2s60_burst_10_downstream_read & ~sys_clk_timer_s1_waits_for_read;

  //sys_clk_timer_s1_writedata mux, which is an e_mux
  assign sys_clk_timer_s1_writedata = std_2s60_burst_10_downstream_writedata;

  //master is always granted when requested
  assign std_2s60_burst_10_downstream_granted_sys_clk_timer_s1 = std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1;

  //std_2s60_burst_10/downstream saved-grant sys_clk_timer/s1, which is an e_assign
  assign std_2s60_burst_10_downstream_saved_grant_sys_clk_timer_s1 = std_2s60_burst_10_downstream_requests_sys_clk_timer_s1;

  //allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  assign sys_clk_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sys_clk_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sys_clk_timer_s1_master_qreq_vector = 1;

  //sys_clk_timer_s1_reset_n assignment, which is an e_assign
  assign sys_clk_timer_s1_reset_n = reset_n;

  assign sys_clk_timer_s1_chipselect = std_2s60_burst_10_downstream_granted_sys_clk_timer_s1;
  //sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  assign sys_clk_timer_s1_firsttransfer = sys_clk_timer_s1_begins_xfer ? sys_clk_timer_s1_unreg_firsttransfer : sys_clk_timer_s1_reg_firsttransfer;

  //sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sys_clk_timer_s1_unreg_firsttransfer = ~(sys_clk_timer_s1_slavearbiterlockenable & sys_clk_timer_s1_any_continuerequest);

  //sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_reg_firsttransfer <= 1'b1;
      else if (sys_clk_timer_s1_begins_xfer)
          sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
    end


  //sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sys_clk_timer_s1_beginbursttransfer_internal = sys_clk_timer_s1_begins_xfer;

  //~sys_clk_timer_s1_write_n assignment, which is an e_mux
  assign sys_clk_timer_s1_write_n = ~(std_2s60_burst_10_downstream_granted_sys_clk_timer_s1 & std_2s60_burst_10_downstream_write);

  //sys_clk_timer_s1_address mux, which is an e_mux
  assign sys_clk_timer_s1_address = std_2s60_burst_10_downstream_nativeaddress;

  //d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sys_clk_timer_s1_end_xfer <= 1;
      else if (1)
          d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end


  //sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign sys_clk_timer_s1_waits_for_read = sys_clk_timer_s1_in_a_read_cycle & sys_clk_timer_s1_begins_xfer;

  //sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign sys_clk_timer_s1_in_a_read_cycle = std_2s60_burst_10_downstream_granted_sys_clk_timer_s1 & std_2s60_burst_10_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sys_clk_timer_s1_in_a_read_cycle;

  //sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign sys_clk_timer_s1_waits_for_write = sys_clk_timer_s1_in_a_write_cycle & 0;

  //sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign sys_clk_timer_s1_in_a_write_cycle = std_2s60_burst_10_downstream_granted_sys_clk_timer_s1 & std_2s60_burst_10_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sys_clk_timer_s1_in_a_write_cycle;

  assign wait_for_sys_clk_timer_s1_counter = 0;
  //assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sys_clk_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_10/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_10_downstream_requests_sys_clk_timer_s1 && (std_2s60_burst_10_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_10/downstream drove 0 on its 'arbitrationshare' port while accessing slave sys_clk_timer/s1", $time);
          $stop;
        end
    end


  //std_2s60_burst_10/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_10_downstream_requests_sys_clk_timer_s1 && (std_2s60_burst_10_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_10/downstream drove 0 on its 'burstcount' port while accessing slave sys_clk_timer/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         reset_n,
                                         std_2s60_burst_14_downstream_address_to_slave,
                                         std_2s60_burst_14_downstream_arbitrationshare,
                                         std_2s60_burst_14_downstream_burstcount,
                                         std_2s60_burst_14_downstream_latency_counter,
                                         std_2s60_burst_14_downstream_nativeaddress,
                                         std_2s60_burst_14_downstream_read,
                                         std_2s60_burst_14_downstream_write,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         d1_sysid_control_slave_end_xfer,
                                         std_2s60_burst_14_downstream_granted_sysid_control_slave,
                                         std_2s60_burst_14_downstream_qualified_request_sysid_control_slave,
                                         std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave,
                                         std_2s60_burst_14_downstream_requests_sysid_control_slave,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa
                                      )
;

  output           d1_sysid_control_slave_end_xfer;
  output           std_2s60_burst_14_downstream_granted_sysid_control_slave;
  output           std_2s60_burst_14_downstream_qualified_request_sysid_control_slave;
  output           std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave;
  output           std_2s60_burst_14_downstream_requests_sysid_control_slave;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  input            clk;
  input            reset_n;
  input   [  2: 0] std_2s60_burst_14_downstream_address_to_slave;
  input   [  3: 0] std_2s60_burst_14_downstream_arbitrationshare;
  input            std_2s60_burst_14_downstream_burstcount;
  input            std_2s60_burst_14_downstream_latency_counter;
  input   [  2: 0] std_2s60_burst_14_downstream_nativeaddress;
  input            std_2s60_burst_14_downstream_read;
  input            std_2s60_burst_14_downstream_write;
  input   [ 31: 0] sysid_control_slave_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             std_2s60_burst_14_downstream_arbiterlock;
  wire             std_2s60_burst_14_downstream_arbiterlock2;
  wire             std_2s60_burst_14_downstream_continuerequest;
  wire             std_2s60_burst_14_downstream_granted_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_qualified_request_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_requests_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_saved_grant_sysid_control_slave;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg     [  3: 0] sysid_control_slave_arb_share_counter;
  wire    [  3: 0] sysid_control_slave_arb_share_counter_next_value;
  wire    [  3: 0] sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else if (1)
          d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((std_2s60_burst_14_downstream_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign std_2s60_burst_14_downstream_requests_sysid_control_slave = ((1) & (std_2s60_burst_14_downstream_read | std_2s60_burst_14_downstream_write)) & std_2s60_burst_14_downstream_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = (std_2s60_burst_14_downstream_granted_sysid_control_slave)? std_2s60_burst_14_downstream_arbitrationshare :
    1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = 0;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = std_2s60_burst_14_downstream_saved_grant_sysid_control_slave;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //std_2s60_burst_14/downstream sysid/control_slave arbiterlock, which is an e_assign
  assign std_2s60_burst_14_downstream_arbiterlock = sysid_control_slave_slavearbiterlockenable & std_2s60_burst_14_downstream_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //std_2s60_burst_14/downstream sysid/control_slave arbiterlock2, which is an e_assign
  assign std_2s60_burst_14_downstream_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & std_2s60_burst_14_downstream_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //std_2s60_burst_14_downstream_continuerequest continued request, which is an e_assign
  assign std_2s60_burst_14_downstream_continuerequest = 1;

  assign std_2s60_burst_14_downstream_qualified_request_sysid_control_slave = std_2s60_burst_14_downstream_requests_sysid_control_slave & ~((std_2s60_burst_14_downstream_read & ((std_2s60_burst_14_downstream_latency_counter != 0))));
  //local readdatavalid std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave, which is an e_mux
  assign std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave = std_2s60_burst_14_downstream_granted_sysid_control_slave & std_2s60_burst_14_downstream_read & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign std_2s60_burst_14_downstream_granted_sysid_control_slave = std_2s60_burst_14_downstream_qualified_request_sysid_control_slave;

  //std_2s60_burst_14/downstream saved-grant sysid/control_slave, which is an e_assign
  assign std_2s60_burst_14_downstream_saved_grant_sysid_control_slave = std_2s60_burst_14_downstream_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = std_2s60_burst_14_downstream_nativeaddress;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else if (1)
          d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = std_2s60_burst_14_downstream_granted_sysid_control_slave & std_2s60_burst_14_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = std_2s60_burst_14_downstream_granted_sysid_control_slave & std_2s60_burst_14_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else if (1)
          enable_nonzero_assertions <= 1'b1;
    end


  //std_2s60_burst_14/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_14_downstream_requests_sysid_control_slave && (std_2s60_burst_14_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_14/downstream drove 0 on its 'arbitrationshare' port while accessing slave sysid/control_slave", $time);
          $stop;
        end
    end


  //std_2s60_burst_14/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (std_2s60_burst_14_downstream_requests_sysid_control_slave && (std_2s60_burst_14_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: std_2s60_burst_14/downstream drove 0 on its 'burstcount' port while accessing slave sysid/control_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60_reset_clk_domain_synch_module (
                                                // inputs:
                                                 clk,
                                                 data_in,
                                                 reset_n,

                                                // outputs:
                                                 data_out
                                              )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else if (1)
          data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else if (1)
          data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module std_2s60 (
                  // 1) global signals:
                   clk,
                   reset_n,

                  // the_ad_buf
                   a2dc_to_the_ad_buf,
                   adclk_to_the_ad_buf,
                   wrclk_to_the_ad_buf,

                  // the_ext_flash_bus_avalon_slave
                   ext_flash_bus_address,
                   ext_flash_bus_data,
                   ext_flash_bus_readn,
                   select_n_to_the_ext_flash,
                   write_n_to_the_ext_flash,

                  // the_ext_ram_bus_avalon_slave
                   be_n_to_the_ext_ram,
                   ext_ram_bus_address,
                   ext_ram_bus_byteenablen,
                   ext_ram_bus_data,
                   ior_n_to_the_lan91c111,
                   iow_n_to_the_lan91c111,
                   irq_from_the_lan91c111,
                   read_n_to_the_ext_ram,
                   reset_to_the_lan91c111,
                   select_n_to_the_ext_ram,
                   write_n_to_the_ext_ram,

                  // the_reconfig_request_pio
                   bidir_port_to_and_from_the_reconfig_request_pio,

                  // the_sdram
                   zs_addr_from_the_sdram,
                   zs_ba_from_the_sdram,
                   zs_cas_n_from_the_sdram,
                   zs_cke_from_the_sdram,
                   zs_cs_n_from_the_sdram,
                   zs_dq_to_and_from_the_sdram,
                   zs_dqm_from_the_sdram,
                   zs_ras_n_from_the_sdram,
                   zs_we_n_from_the_sdram
                )
;

  output  [  3: 0] be_n_to_the_ext_ram;
  inout            bidir_port_to_and_from_the_reconfig_request_pio;
  output  [ 23: 0] ext_flash_bus_address;
  inout   [  7: 0] ext_flash_bus_data;
  output           ext_flash_bus_readn;
  output  [ 19: 0] ext_ram_bus_address;
  output  [  3: 0] ext_ram_bus_byteenablen;
  inout   [ 31: 0] ext_ram_bus_data;
  output           ior_n_to_the_lan91c111;
  output           iow_n_to_the_lan91c111;
  output           read_n_to_the_ext_ram;
  output           reset_to_the_lan91c111;
  output           select_n_to_the_ext_flash;
  output           select_n_to_the_ext_ram;
  output           write_n_to_the_ext_flash;
  output           write_n_to_the_ext_ram;
  output  [ 11: 0] zs_addr_from_the_sdram;
  output  [  1: 0] zs_ba_from_the_sdram;
  output           zs_cas_n_from_the_sdram;
  output           zs_cke_from_the_sdram;
  output           zs_cs_n_from_the_sdram;
  inout   [ 31: 0] zs_dq_to_and_from_the_sdram;
  output  [  3: 0] zs_dqm_from_the_sdram;
  output           zs_ras_n_from_the_sdram;
  output           zs_we_n_from_the_sdram;
  input   [ 11: 0] a2dc_to_the_ad_buf;
  input            adclk_to_the_ad_buf;
  input            clk;
  input            irq_from_the_lan91c111;
  input            reset_n;
  input            wrclk_to_the_ad_buf;

  wire    [ 11: 0] ad_buf_s1_address;
  wire             ad_buf_s1_chipselect_n;
  wire             ad_buf_s1_read;
  wire    [ 31: 0] ad_buf_s1_readdata;
  wire    [ 31: 0] ad_buf_s1_readdata_from_sa;
  wire             ad_buf_s1_reset_n;
  wire             ad_buf_s1_waitrequest;
  wire             ad_buf_s1_waitrequest_from_sa;
  wire    [  3: 0] be_n_to_the_ext_ram;
  wire             bidir_port_to_and_from_the_reconfig_request_pio;
  wire             clk_reset_n;
  wire    [ 25: 0] cpu_data_master_address;
  wire    [ 25: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_burstcount;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire             cpu_data_master_byteenable_std_2s60_burst_3_upstream;
  wire    [  1: 0] cpu_data_master_dbs_address;
  wire    [  7: 0] cpu_data_master_dbs_write_8;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_std_2s60_burst_10_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_11_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_12_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_13_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_14_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_16_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_17_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_1_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_3_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_5_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_7_upstream;
  wire             cpu_data_master_granted_std_2s60_burst_9_upstream;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_std_2s60_burst_10_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_11_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_12_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_13_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_14_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_16_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_17_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_1_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_3_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_5_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_7_upstream;
  wire             cpu_data_master_qualified_request_std_2s60_burst_9_upstream;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_10_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_11_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_12_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_13_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_14_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_16_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_17_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_1_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_3_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_5_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_7_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_9_upstream;
  wire             cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_std_2s60_burst_10_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_11_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_12_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_13_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_14_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_16_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_17_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_1_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_3_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_5_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_7_upstream;
  wire             cpu_data_master_requests_std_2s60_burst_9_upstream;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 25: 0] cpu_instruction_master_address;
  wire    [ 25: 0] cpu_instruction_master_address_to_slave;
  wire    [  3: 0] cpu_instruction_master_burstcount;
  wire    [  1: 0] cpu_instruction_master_dbs_address;
  wire             cpu_instruction_master_granted_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_granted_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_std_2s60_burst_0_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_15_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_18_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_2_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_4_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_6_upstream;
  wire             cpu_instruction_master_requests_std_2s60_burst_8_upstream;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire             d1_ad_buf_s1_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_ext_flash_bus_avalon_slave_end_xfer;
  wire             d1_ext_ram_bus_avalon_slave_end_xfer;
  wire             d1_high_res_timer_s1_end_xfer;
  wire             d1_irq_from_the_lan91c111;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_onchip_ram_64_kbytes_s1_end_xfer;
  wire             d1_reconfig_request_pio_s1_end_xfer;
  wire             d1_sdram_s1_end_xfer;
  wire             d1_std_2s60_burst_0_upstream_end_xfer;
  wire             d1_std_2s60_burst_10_upstream_end_xfer;
  wire             d1_std_2s60_burst_11_upstream_end_xfer;
  wire             d1_std_2s60_burst_12_upstream_end_xfer;
  wire             d1_std_2s60_burst_13_upstream_end_xfer;
  wire             d1_std_2s60_burst_14_upstream_end_xfer;
  wire             d1_std_2s60_burst_15_upstream_end_xfer;
  wire             d1_std_2s60_burst_16_upstream_end_xfer;
  wire             d1_std_2s60_burst_17_upstream_end_xfer;
  wire             d1_std_2s60_burst_18_upstream_end_xfer;
  wire             d1_std_2s60_burst_1_upstream_end_xfer;
  wire             d1_std_2s60_burst_2_upstream_end_xfer;
  wire             d1_std_2s60_burst_3_upstream_end_xfer;
  wire             d1_std_2s60_burst_4_upstream_end_xfer;
  wire             d1_std_2s60_burst_5_upstream_end_xfer;
  wire             d1_std_2s60_burst_6_upstream_end_xfer;
  wire             d1_std_2s60_burst_7_upstream_end_xfer;
  wire             d1_std_2s60_burst_8_upstream_end_xfer;
  wire             d1_std_2s60_burst_9_upstream_end_xfer;
  wire             d1_sys_clk_timer_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire    [ 23: 0] ext_flash_bus_address;
  wire    [  7: 0] ext_flash_bus_data;
  wire             ext_flash_bus_readn;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire    [ 19: 0] ext_ram_bus_address;
  wire    [  3: 0] ext_ram_bus_byteenablen;
  wire    [ 31: 0] ext_ram_bus_data;
  wire             ext_ram_s1_wait_counter_eq_0;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_irq;
  wire             high_res_timer_s1_irq_from_sa;
  wire    [ 15: 0] high_res_timer_s1_readdata;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  wire             high_res_timer_s1_reset_n;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire    [  7: 0] incoming_ext_flash_bus_data_with_Xs_converted_to_0;
  wire    [ 31: 0] incoming_ext_ram_bus_data;
  wire             ior_n_to_the_lan91c111;
  wire             iow_n_to_the_lan91c111;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             lan91c111_s1_wait_counter_eq_0;
  wire    [ 13: 0] onchip_ram_64_kbytes_s1_address;
  wire    [  3: 0] onchip_ram_64_kbytes_s1_byteenable;
  wire             onchip_ram_64_kbytes_s1_chipselect;
  wire             onchip_ram_64_kbytes_s1_clken;
  wire    [ 31: 0] onchip_ram_64_kbytes_s1_readdata;
  wire    [ 31: 0] onchip_ram_64_kbytes_s1_readdata_from_sa;
  wire             onchip_ram_64_kbytes_s1_write;
  wire    [ 31: 0] onchip_ram_64_kbytes_s1_writedata;
  wire             read_n_to_the_ext_ram;
  wire    [  1: 0] reconfig_request_pio_s1_address;
  wire             reconfig_request_pio_s1_chipselect;
  wire             reconfig_request_pio_s1_readdata;
  wire             reconfig_request_pio_s1_readdata_from_sa;
  wire             reconfig_request_pio_s1_reset_n;
  wire             reconfig_request_pio_s1_write_n;
  wire             reconfig_request_pio_s1_writedata;
  wire             reset_n_sources;
  wire             reset_to_the_lan91c111;
  wire    [ 21: 0] sdram_s1_address;
  wire    [  3: 0] sdram_s1_byteenable_n;
  wire             sdram_s1_chipselect;
  wire             sdram_s1_read_n;
  wire    [ 31: 0] sdram_s1_readdata;
  wire    [ 31: 0] sdram_s1_readdata_from_sa;
  wire             sdram_s1_readdatavalid;
  wire             sdram_s1_reset_n;
  wire             sdram_s1_waitrequest;
  wire             sdram_s1_waitrequest_from_sa;
  wire             sdram_s1_write_n;
  wire    [ 31: 0] sdram_s1_writedata;
  wire             select_n_to_the_ext_flash;
  wire             select_n_to_the_ext_ram;
  wire    [ 10: 0] std_2s60_burst_0_downstream_address;
  wire    [ 10: 0] std_2s60_burst_0_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_0_downstream_arbitrationshare;
  wire             std_2s60_burst_0_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_0_downstream_byteenable;
  wire             std_2s60_burst_0_downstream_debugaccess;
  wire             std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_latency_counter;
  wire    [ 10: 0] std_2s60_burst_0_downstream_nativeaddress;
  wire             std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_read;
  wire             std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module;
  wire    [ 31: 0] std_2s60_burst_0_downstream_readdata;
  wire             std_2s60_burst_0_downstream_readdatavalid;
  wire             std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module;
  wire             std_2s60_burst_0_downstream_reset_n;
  wire             std_2s60_burst_0_downstream_waitrequest;
  wire             std_2s60_burst_0_downstream_write;
  wire    [ 31: 0] std_2s60_burst_0_downstream_writedata;
  wire    [ 10: 0] std_2s60_burst_0_upstream_address;
  wire    [ 12: 0] std_2s60_burst_0_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_0_upstream_byteenable;
  wire             std_2s60_burst_0_upstream_debugaccess;
  wire             std_2s60_burst_0_upstream_read;
  wire    [ 31: 0] std_2s60_burst_0_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_0_upstream_readdata_from_sa;
  wire             std_2s60_burst_0_upstream_readdatavalid;
  wire             std_2s60_burst_0_upstream_waitrequest;
  wire             std_2s60_burst_0_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_0_upstream_write;
  wire    [ 31: 0] std_2s60_burst_0_upstream_writedata;
  wire    [  3: 0] std_2s60_burst_10_downstream_address;
  wire    [  3: 0] std_2s60_burst_10_downstream_address_to_slave;
  wire    [  4: 0] std_2s60_burst_10_downstream_arbitrationshare;
  wire             std_2s60_burst_10_downstream_burstcount;
  wire    [  1: 0] std_2s60_burst_10_downstream_byteenable;
  wire             std_2s60_burst_10_downstream_debugaccess;
  wire             std_2s60_burst_10_downstream_granted_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_latency_counter;
  wire    [  3: 0] std_2s60_burst_10_downstream_nativeaddress;
  wire             std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_read;
  wire             std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1;
  wire    [ 15: 0] std_2s60_burst_10_downstream_readdata;
  wire             std_2s60_burst_10_downstream_readdatavalid;
  wire             std_2s60_burst_10_downstream_requests_sys_clk_timer_s1;
  wire             std_2s60_burst_10_downstream_reset_n;
  wire             std_2s60_burst_10_downstream_waitrequest;
  wire             std_2s60_burst_10_downstream_write;
  wire    [ 15: 0] std_2s60_burst_10_downstream_writedata;
  wire    [  3: 0] std_2s60_burst_10_upstream_address;
  wire    [  3: 0] std_2s60_burst_10_upstream_burstcount;
  wire    [  4: 0] std_2s60_burst_10_upstream_byteaddress;
  wire    [  1: 0] std_2s60_burst_10_upstream_byteenable;
  wire             std_2s60_burst_10_upstream_debugaccess;
  wire             std_2s60_burst_10_upstream_read;
  wire    [ 15: 0] std_2s60_burst_10_upstream_readdata;
  wire    [ 15: 0] std_2s60_burst_10_upstream_readdata_from_sa;
  wire             std_2s60_burst_10_upstream_readdatavalid;
  wire             std_2s60_burst_10_upstream_waitrequest;
  wire             std_2s60_burst_10_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_10_upstream_write;
  wire    [ 15: 0] std_2s60_burst_10_upstream_writedata;
  wire    [  2: 0] std_2s60_burst_11_downstream_address;
  wire    [  2: 0] std_2s60_burst_11_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_11_downstream_arbitrationshare;
  wire             std_2s60_burst_11_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_11_downstream_byteenable;
  wire             std_2s60_burst_11_downstream_debugaccess;
  wire             std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_latency_counter;
  wire    [  2: 0] std_2s60_burst_11_downstream_nativeaddress;
  wire             std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_read;
  wire             std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire    [ 31: 0] std_2s60_burst_11_downstream_readdata;
  wire             std_2s60_burst_11_downstream_readdatavalid;
  wire             std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave;
  wire             std_2s60_burst_11_downstream_reset_n;
  wire             std_2s60_burst_11_downstream_waitrequest;
  wire             std_2s60_burst_11_downstream_write;
  wire    [ 31: 0] std_2s60_burst_11_downstream_writedata;
  wire    [  2: 0] std_2s60_burst_11_upstream_address;
  wire    [  3: 0] std_2s60_burst_11_upstream_burstcount;
  wire    [  4: 0] std_2s60_burst_11_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_11_upstream_byteenable;
  wire             std_2s60_burst_11_upstream_debugaccess;
  wire             std_2s60_burst_11_upstream_read;
  wire    [ 31: 0] std_2s60_burst_11_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_11_upstream_readdata_from_sa;
  wire             std_2s60_burst_11_upstream_readdatavalid;
  wire             std_2s60_burst_11_upstream_waitrequest;
  wire             std_2s60_burst_11_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_11_upstream_write;
  wire    [ 31: 0] std_2s60_burst_11_upstream_writedata;
  wire    [  3: 0] std_2s60_burst_12_downstream_address;
  wire    [  3: 0] std_2s60_burst_12_downstream_address_to_slave;
  wire    [  4: 0] std_2s60_burst_12_downstream_arbitrationshare;
  wire             std_2s60_burst_12_downstream_burstcount;
  wire    [  1: 0] std_2s60_burst_12_downstream_byteenable;
  wire             std_2s60_burst_12_downstream_debugaccess;
  wire             std_2s60_burst_12_downstream_granted_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_latency_counter;
  wire    [  3: 0] std_2s60_burst_12_downstream_nativeaddress;
  wire             std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_read;
  wire             std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1;
  wire    [ 15: 0] std_2s60_burst_12_downstream_readdata;
  wire             std_2s60_burst_12_downstream_readdatavalid;
  wire             std_2s60_burst_12_downstream_requests_high_res_timer_s1;
  wire             std_2s60_burst_12_downstream_reset_n;
  wire             std_2s60_burst_12_downstream_waitrequest;
  wire             std_2s60_burst_12_downstream_write;
  wire    [ 15: 0] std_2s60_burst_12_downstream_writedata;
  wire    [  3: 0] std_2s60_burst_12_upstream_address;
  wire    [  3: 0] std_2s60_burst_12_upstream_burstcount;
  wire    [  4: 0] std_2s60_burst_12_upstream_byteaddress;
  wire    [  1: 0] std_2s60_burst_12_upstream_byteenable;
  wire             std_2s60_burst_12_upstream_debugaccess;
  wire             std_2s60_burst_12_upstream_read;
  wire    [ 15: 0] std_2s60_burst_12_upstream_readdata;
  wire    [ 15: 0] std_2s60_burst_12_upstream_readdata_from_sa;
  wire             std_2s60_burst_12_upstream_readdatavalid;
  wire             std_2s60_burst_12_upstream_waitrequest;
  wire             std_2s60_burst_12_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_12_upstream_write;
  wire    [ 15: 0] std_2s60_burst_12_upstream_writedata;
  wire    [  1: 0] std_2s60_burst_13_downstream_address;
  wire    [  1: 0] std_2s60_burst_13_downstream_address_to_slave;
  wire    [  5: 0] std_2s60_burst_13_downstream_arbitrationshare;
  wire             std_2s60_burst_13_downstream_burstcount;
  wire             std_2s60_burst_13_downstream_byteenable;
  wire             std_2s60_burst_13_downstream_debugaccess;
  wire             std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_latency_counter;
  wire    [  1: 0] std_2s60_burst_13_downstream_nativeaddress;
  wire             std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_read;
  wire             std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1;
  wire    [  7: 0] std_2s60_burst_13_downstream_readdata;
  wire             std_2s60_burst_13_downstream_readdatavalid;
  wire             std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1;
  wire             std_2s60_burst_13_downstream_reset_n;
  wire             std_2s60_burst_13_downstream_waitrequest;
  wire             std_2s60_burst_13_downstream_write;
  wire    [  7: 0] std_2s60_burst_13_downstream_writedata;
  wire    [  1: 0] std_2s60_burst_13_upstream_address;
  wire    [  3: 0] std_2s60_burst_13_upstream_burstcount;
  wire    [  1: 0] std_2s60_burst_13_upstream_byteaddress;
  wire             std_2s60_burst_13_upstream_byteenable;
  wire             std_2s60_burst_13_upstream_debugaccess;
  wire             std_2s60_burst_13_upstream_read;
  wire    [  7: 0] std_2s60_burst_13_upstream_readdata;
  wire    [  7: 0] std_2s60_burst_13_upstream_readdata_from_sa;
  wire             std_2s60_burst_13_upstream_readdatavalid;
  wire             std_2s60_burst_13_upstream_waitrequest;
  wire             std_2s60_burst_13_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_13_upstream_write;
  wire    [  7: 0] std_2s60_burst_13_upstream_writedata;
  wire    [  2: 0] std_2s60_burst_14_downstream_address;
  wire    [  2: 0] std_2s60_burst_14_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_14_downstream_arbitrationshare;
  wire             std_2s60_burst_14_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_14_downstream_byteenable;
  wire             std_2s60_burst_14_downstream_debugaccess;
  wire             std_2s60_burst_14_downstream_granted_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_latency_counter;
  wire    [  2: 0] std_2s60_burst_14_downstream_nativeaddress;
  wire             std_2s60_burst_14_downstream_qualified_request_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_read;
  wire             std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave;
  wire    [ 31: 0] std_2s60_burst_14_downstream_readdata;
  wire             std_2s60_burst_14_downstream_readdatavalid;
  wire             std_2s60_burst_14_downstream_requests_sysid_control_slave;
  wire             std_2s60_burst_14_downstream_reset_n;
  wire             std_2s60_burst_14_downstream_waitrequest;
  wire             std_2s60_burst_14_downstream_write;
  wire    [ 31: 0] std_2s60_burst_14_downstream_writedata;
  wire    [  2: 0] std_2s60_burst_14_upstream_address;
  wire    [  3: 0] std_2s60_burst_14_upstream_burstcount;
  wire    [  4: 0] std_2s60_burst_14_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_14_upstream_byteenable;
  wire             std_2s60_burst_14_upstream_debugaccess;
  wire             std_2s60_burst_14_upstream_read;
  wire    [ 31: 0] std_2s60_burst_14_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_14_upstream_readdata_from_sa;
  wire             std_2s60_burst_14_upstream_readdatavalid;
  wire             std_2s60_burst_14_upstream_waitrequest;
  wire             std_2s60_burst_14_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_14_upstream_write;
  wire    [ 31: 0] std_2s60_burst_14_upstream_writedata;
  wire    [ 23: 0] std_2s60_burst_15_downstream_address;
  wire    [ 23: 0] std_2s60_burst_15_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_15_downstream_arbitrationshare;
  wire             std_2s60_burst_15_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_15_downstream_byteenable;
  wire             std_2s60_burst_15_downstream_debugaccess;
  wire             std_2s60_burst_15_downstream_granted_sdram_s1;
  wire             std_2s60_burst_15_downstream_latency_counter;
  wire    [ 23: 0] std_2s60_burst_15_downstream_nativeaddress;
  wire             std_2s60_burst_15_downstream_qualified_request_sdram_s1;
  wire             std_2s60_burst_15_downstream_read;
  wire             std_2s60_burst_15_downstream_read_data_valid_sdram_s1;
  wire             std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register;
  wire    [ 31: 0] std_2s60_burst_15_downstream_readdata;
  wire             std_2s60_burst_15_downstream_readdatavalid;
  wire             std_2s60_burst_15_downstream_requests_sdram_s1;
  wire             std_2s60_burst_15_downstream_reset_n;
  wire             std_2s60_burst_15_downstream_waitrequest;
  wire             std_2s60_burst_15_downstream_write;
  wire    [ 31: 0] std_2s60_burst_15_downstream_writedata;
  wire    [ 23: 0] std_2s60_burst_15_upstream_address;
  wire    [ 25: 0] std_2s60_burst_15_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_15_upstream_byteenable;
  wire             std_2s60_burst_15_upstream_debugaccess;
  wire             std_2s60_burst_15_upstream_read;
  wire    [ 31: 0] std_2s60_burst_15_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_15_upstream_readdata_from_sa;
  wire             std_2s60_burst_15_upstream_readdatavalid;
  wire             std_2s60_burst_15_upstream_waitrequest;
  wire             std_2s60_burst_15_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_15_upstream_write;
  wire    [ 31: 0] std_2s60_burst_15_upstream_writedata;
  wire    [ 23: 0] std_2s60_burst_16_downstream_address;
  wire    [ 23: 0] std_2s60_burst_16_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_16_downstream_arbitrationshare;
  wire             std_2s60_burst_16_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_16_downstream_byteenable;
  wire             std_2s60_burst_16_downstream_debugaccess;
  wire             std_2s60_burst_16_downstream_granted_sdram_s1;
  wire             std_2s60_burst_16_downstream_latency_counter;
  wire    [ 23: 0] std_2s60_burst_16_downstream_nativeaddress;
  wire             std_2s60_burst_16_downstream_qualified_request_sdram_s1;
  wire             std_2s60_burst_16_downstream_read;
  wire             std_2s60_burst_16_downstream_read_data_valid_sdram_s1;
  wire             std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register;
  wire    [ 31: 0] std_2s60_burst_16_downstream_readdata;
  wire             std_2s60_burst_16_downstream_readdatavalid;
  wire             std_2s60_burst_16_downstream_requests_sdram_s1;
  wire             std_2s60_burst_16_downstream_reset_n;
  wire             std_2s60_burst_16_downstream_waitrequest;
  wire             std_2s60_burst_16_downstream_write;
  wire    [ 31: 0] std_2s60_burst_16_downstream_writedata;
  wire    [ 23: 0] std_2s60_burst_16_upstream_address;
  wire    [  3: 0] std_2s60_burst_16_upstream_burstcount;
  wire    [ 25: 0] std_2s60_burst_16_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_16_upstream_byteenable;
  wire             std_2s60_burst_16_upstream_debugaccess;
  wire             std_2s60_burst_16_upstream_read;
  wire    [ 31: 0] std_2s60_burst_16_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_16_upstream_readdata_from_sa;
  wire             std_2s60_burst_16_upstream_readdatavalid;
  wire             std_2s60_burst_16_upstream_waitrequest;
  wire             std_2s60_burst_16_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_16_upstream_write;
  wire    [ 31: 0] std_2s60_burst_16_upstream_writedata;
  wire    [ 13: 0] std_2s60_burst_17_downstream_address;
  wire    [ 13: 0] std_2s60_burst_17_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_17_downstream_arbitrationshare;
  wire             std_2s60_burst_17_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_17_downstream_byteenable;
  wire             std_2s60_burst_17_downstream_debugaccess;
  wire             std_2s60_burst_17_downstream_granted_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_latency_counter;
  wire    [ 13: 0] std_2s60_burst_17_downstream_nativeaddress;
  wire             std_2s60_burst_17_downstream_qualified_request_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_read;
  wire             std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1;
  wire    [ 31: 0] std_2s60_burst_17_downstream_readdata;
  wire             std_2s60_burst_17_downstream_readdatavalid;
  wire             std_2s60_burst_17_downstream_requests_ad_buf_s1;
  wire             std_2s60_burst_17_downstream_reset_n;
  wire             std_2s60_burst_17_downstream_waitrequest;
  wire             std_2s60_burst_17_downstream_write;
  wire    [ 31: 0] std_2s60_burst_17_downstream_writedata;
  wire    [ 13: 0] std_2s60_burst_17_upstream_address;
  wire    [  3: 0] std_2s60_burst_17_upstream_burstcount;
  wire    [ 15: 0] std_2s60_burst_17_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_17_upstream_byteenable;
  wire             std_2s60_burst_17_upstream_debugaccess;
  wire             std_2s60_burst_17_upstream_read;
  wire    [ 31: 0] std_2s60_burst_17_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_17_upstream_readdata_from_sa;
  wire             std_2s60_burst_17_upstream_readdatavalid;
  wire             std_2s60_burst_17_upstream_waitrequest;
  wire             std_2s60_burst_17_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_17_upstream_write;
  wire    [ 31: 0] std_2s60_burst_17_upstream_writedata;
  wire    [ 13: 0] std_2s60_burst_18_downstream_address;
  wire    [ 13: 0] std_2s60_burst_18_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_18_downstream_arbitrationshare;
  wire             std_2s60_burst_18_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_18_downstream_byteenable;
  wire             std_2s60_burst_18_downstream_debugaccess;
  wire             std_2s60_burst_18_downstream_granted_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_latency_counter;
  wire    [ 13: 0] std_2s60_burst_18_downstream_nativeaddress;
  wire             std_2s60_burst_18_downstream_qualified_request_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_read;
  wire             std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1;
  wire    [ 31: 0] std_2s60_burst_18_downstream_readdata;
  wire             std_2s60_burst_18_downstream_readdatavalid;
  wire             std_2s60_burst_18_downstream_requests_ad_buf_s1;
  wire             std_2s60_burst_18_downstream_reset_n;
  wire             std_2s60_burst_18_downstream_waitrequest;
  wire             std_2s60_burst_18_downstream_write;
  wire    [ 31: 0] std_2s60_burst_18_downstream_writedata;
  wire    [ 13: 0] std_2s60_burst_18_upstream_address;
  wire    [ 15: 0] std_2s60_burst_18_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_18_upstream_byteenable;
  wire             std_2s60_burst_18_upstream_debugaccess;
  wire             std_2s60_burst_18_upstream_read;
  wire    [ 31: 0] std_2s60_burst_18_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_18_upstream_readdata_from_sa;
  wire             std_2s60_burst_18_upstream_readdatavalid;
  wire             std_2s60_burst_18_upstream_waitrequest;
  wire             std_2s60_burst_18_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_18_upstream_write;
  wire    [ 31: 0] std_2s60_burst_18_upstream_writedata;
  wire    [ 10: 0] std_2s60_burst_1_downstream_address;
  wire    [ 10: 0] std_2s60_burst_1_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_1_downstream_arbitrationshare;
  wire             std_2s60_burst_1_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_1_downstream_byteenable;
  wire             std_2s60_burst_1_downstream_debugaccess;
  wire             std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_latency_counter;
  wire    [ 10: 0] std_2s60_burst_1_downstream_nativeaddress;
  wire             std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_read;
  wire             std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module;
  wire    [ 31: 0] std_2s60_burst_1_downstream_readdata;
  wire             std_2s60_burst_1_downstream_readdatavalid;
  wire             std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module;
  wire             std_2s60_burst_1_downstream_reset_n;
  wire             std_2s60_burst_1_downstream_waitrequest;
  wire             std_2s60_burst_1_downstream_write;
  wire    [ 31: 0] std_2s60_burst_1_downstream_writedata;
  wire    [ 10: 0] std_2s60_burst_1_upstream_address;
  wire    [  3: 0] std_2s60_burst_1_upstream_burstcount;
  wire    [ 12: 0] std_2s60_burst_1_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_1_upstream_byteenable;
  wire             std_2s60_burst_1_upstream_debugaccess;
  wire             std_2s60_burst_1_upstream_read;
  wire    [ 31: 0] std_2s60_burst_1_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_1_upstream_readdata_from_sa;
  wire             std_2s60_burst_1_upstream_readdatavalid;
  wire             std_2s60_burst_1_upstream_waitrequest;
  wire             std_2s60_burst_1_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_1_upstream_write;
  wire    [ 31: 0] std_2s60_burst_1_upstream_writedata;
  wire    [ 23: 0] std_2s60_burst_2_downstream_address;
  wire    [ 23: 0] std_2s60_burst_2_downstream_address_to_slave;
  wire    [  5: 0] std_2s60_burst_2_downstream_arbitrationshare;
  wire             std_2s60_burst_2_downstream_burstcount;
  wire             std_2s60_burst_2_downstream_byteenable;
  wire             std_2s60_burst_2_downstream_debugaccess;
  wire             std_2s60_burst_2_downstream_granted_ext_flash_s1;
  wire    [  1: 0] std_2s60_burst_2_downstream_latency_counter;
  wire    [ 23: 0] std_2s60_burst_2_downstream_nativeaddress;
  wire             std_2s60_burst_2_downstream_qualified_request_ext_flash_s1;
  wire             std_2s60_burst_2_downstream_read;
  wire             std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1;
  wire    [  7: 0] std_2s60_burst_2_downstream_readdata;
  wire             std_2s60_burst_2_downstream_readdatavalid;
  wire             std_2s60_burst_2_downstream_requests_ext_flash_s1;
  wire             std_2s60_burst_2_downstream_reset_n;
  wire             std_2s60_burst_2_downstream_waitrequest;
  wire             std_2s60_burst_2_downstream_write;
  wire    [  7: 0] std_2s60_burst_2_downstream_writedata;
  wire    [ 23: 0] std_2s60_burst_2_upstream_address;
  wire    [ 23: 0] std_2s60_burst_2_upstream_byteaddress;
  wire             std_2s60_burst_2_upstream_byteenable;
  wire             std_2s60_burst_2_upstream_debugaccess;
  wire             std_2s60_burst_2_upstream_read;
  wire    [  7: 0] std_2s60_burst_2_upstream_readdata;
  wire    [  7: 0] std_2s60_burst_2_upstream_readdata_from_sa;
  wire             std_2s60_burst_2_upstream_readdatavalid;
  wire             std_2s60_burst_2_upstream_waitrequest;
  wire             std_2s60_burst_2_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_2_upstream_write;
  wire    [  7: 0] std_2s60_burst_2_upstream_writedata;
  wire    [ 23: 0] std_2s60_burst_3_downstream_address;
  wire    [ 23: 0] std_2s60_burst_3_downstream_address_to_slave;
  wire    [  5: 0] std_2s60_burst_3_downstream_arbitrationshare;
  wire             std_2s60_burst_3_downstream_burstcount;
  wire             std_2s60_burst_3_downstream_byteenable;
  wire             std_2s60_burst_3_downstream_debugaccess;
  wire             std_2s60_burst_3_downstream_granted_ext_flash_s1;
  wire    [  1: 0] std_2s60_burst_3_downstream_latency_counter;
  wire    [ 23: 0] std_2s60_burst_3_downstream_nativeaddress;
  wire             std_2s60_burst_3_downstream_qualified_request_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_read;
  wire             std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1;
  wire    [  7: 0] std_2s60_burst_3_downstream_readdata;
  wire             std_2s60_burst_3_downstream_readdatavalid;
  wire             std_2s60_burst_3_downstream_requests_ext_flash_s1;
  wire             std_2s60_burst_3_downstream_reset_n;
  wire             std_2s60_burst_3_downstream_waitrequest;
  wire             std_2s60_burst_3_downstream_write;
  wire    [  7: 0] std_2s60_burst_3_downstream_writedata;
  wire    [ 23: 0] std_2s60_burst_3_upstream_address;
  wire    [  3: 0] std_2s60_burst_3_upstream_burstcount;
  wire    [ 23: 0] std_2s60_burst_3_upstream_byteaddress;
  wire             std_2s60_burst_3_upstream_byteenable;
  wire             std_2s60_burst_3_upstream_debugaccess;
  wire             std_2s60_burst_3_upstream_read;
  wire    [  7: 0] std_2s60_burst_3_upstream_readdata;
  wire    [  7: 0] std_2s60_burst_3_upstream_readdata_from_sa;
  wire             std_2s60_burst_3_upstream_readdatavalid;
  wire             std_2s60_burst_3_upstream_waitrequest;
  wire             std_2s60_burst_3_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_3_upstream_write;
  wire    [  7: 0] std_2s60_burst_3_upstream_writedata;
  wire    [ 19: 0] std_2s60_burst_4_downstream_address;
  wire    [ 19: 0] std_2s60_burst_4_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_4_downstream_arbitrationshare;
  wire             std_2s60_burst_4_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_4_downstream_byteenable;
  wire             std_2s60_burst_4_downstream_debugaccess;
  wire             std_2s60_burst_4_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_granted_lan91c111_s1;
  wire    [  1: 0] std_2s60_burst_4_downstream_latency_counter;
  wire    [ 19: 0] std_2s60_burst_4_downstream_nativeaddress;
  wire             std_2s60_burst_4_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_4_downstream_read;
  wire             std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1;
  wire    [ 31: 0] std_2s60_burst_4_downstream_readdata;
  wire             std_2s60_burst_4_downstream_readdatavalid;
  wire             std_2s60_burst_4_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_4_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_4_downstream_reset_n;
  wire             std_2s60_burst_4_downstream_waitrequest;
  wire             std_2s60_burst_4_downstream_write;
  wire    [ 31: 0] std_2s60_burst_4_downstream_writedata;
  wire    [ 19: 0] std_2s60_burst_4_upstream_address;
  wire    [ 21: 0] std_2s60_burst_4_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_4_upstream_byteenable;
  wire             std_2s60_burst_4_upstream_debugaccess;
  wire             std_2s60_burst_4_upstream_read;
  wire    [ 31: 0] std_2s60_burst_4_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_4_upstream_readdata_from_sa;
  wire             std_2s60_burst_4_upstream_readdatavalid;
  wire             std_2s60_burst_4_upstream_waitrequest;
  wire             std_2s60_burst_4_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_4_upstream_write;
  wire    [ 31: 0] std_2s60_burst_4_upstream_writedata;
  wire    [ 19: 0] std_2s60_burst_5_downstream_address;
  wire    [ 19: 0] std_2s60_burst_5_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_5_downstream_arbitrationshare;
  wire             std_2s60_burst_5_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_5_downstream_byteenable;
  wire             std_2s60_burst_5_downstream_debugaccess;
  wire             std_2s60_burst_5_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_granted_lan91c111_s1;
  wire    [  1: 0] std_2s60_burst_5_downstream_latency_counter;
  wire    [ 19: 0] std_2s60_burst_5_downstream_nativeaddress;
  wire             std_2s60_burst_5_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_read;
  wire             std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1;
  wire    [ 31: 0] std_2s60_burst_5_downstream_readdata;
  wire             std_2s60_burst_5_downstream_readdatavalid;
  wire             std_2s60_burst_5_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_5_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_5_downstream_reset_n;
  wire             std_2s60_burst_5_downstream_waitrequest;
  wire             std_2s60_burst_5_downstream_write;
  wire    [ 31: 0] std_2s60_burst_5_downstream_writedata;
  wire    [ 19: 0] std_2s60_burst_5_upstream_address;
  wire    [  3: 0] std_2s60_burst_5_upstream_burstcount;
  wire    [ 21: 0] std_2s60_burst_5_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_5_upstream_byteenable;
  wire             std_2s60_burst_5_upstream_debugaccess;
  wire             std_2s60_burst_5_upstream_read;
  wire    [ 31: 0] std_2s60_burst_5_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_5_upstream_readdata_from_sa;
  wire             std_2s60_burst_5_upstream_readdatavalid;
  wire             std_2s60_burst_5_upstream_waitrequest;
  wire             std_2s60_burst_5_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_5_upstream_write;
  wire    [ 31: 0] std_2s60_burst_5_upstream_writedata;
  wire    [ 15: 0] std_2s60_burst_6_downstream_address;
  wire    [ 15: 0] std_2s60_burst_6_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_6_downstream_arbitrationshare;
  wire             std_2s60_burst_6_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_6_downstream_byteenable;
  wire             std_2s60_burst_6_downstream_debugaccess;
  wire             std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_latency_counter;
  wire    [ 15: 0] std_2s60_burst_6_downstream_nativeaddress;
  wire             std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_read;
  wire             std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  wire    [ 31: 0] std_2s60_burst_6_downstream_readdata;
  wire             std_2s60_burst_6_downstream_readdatavalid;
  wire             std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_6_downstream_reset_n;
  wire             std_2s60_burst_6_downstream_waitrequest;
  wire             std_2s60_burst_6_downstream_write;
  wire    [ 31: 0] std_2s60_burst_6_downstream_writedata;
  wire    [ 15: 0] std_2s60_burst_6_upstream_address;
  wire    [ 17: 0] std_2s60_burst_6_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_6_upstream_byteenable;
  wire             std_2s60_burst_6_upstream_debugaccess;
  wire             std_2s60_burst_6_upstream_read;
  wire    [ 31: 0] std_2s60_burst_6_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_6_upstream_readdata_from_sa;
  wire             std_2s60_burst_6_upstream_readdatavalid;
  wire             std_2s60_burst_6_upstream_waitrequest;
  wire             std_2s60_burst_6_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_6_upstream_write;
  wire    [ 31: 0] std_2s60_burst_6_upstream_writedata;
  wire    [ 15: 0] std_2s60_burst_7_downstream_address;
  wire    [ 15: 0] std_2s60_burst_7_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_7_downstream_arbitrationshare;
  wire             std_2s60_burst_7_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_7_downstream_byteenable;
  wire             std_2s60_burst_7_downstream_debugaccess;
  wire             std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_latency_counter;
  wire    [ 15: 0] std_2s60_burst_7_downstream_nativeaddress;
  wire             std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_read;
  wire             std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1;
  wire    [ 31: 0] std_2s60_burst_7_downstream_readdata;
  wire             std_2s60_burst_7_downstream_readdatavalid;
  wire             std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1;
  wire             std_2s60_burst_7_downstream_reset_n;
  wire             std_2s60_burst_7_downstream_waitrequest;
  wire             std_2s60_burst_7_downstream_write;
  wire    [ 31: 0] std_2s60_burst_7_downstream_writedata;
  wire    [ 15: 0] std_2s60_burst_7_upstream_address;
  wire    [  3: 0] std_2s60_burst_7_upstream_burstcount;
  wire    [ 17: 0] std_2s60_burst_7_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_7_upstream_byteenable;
  wire             std_2s60_burst_7_upstream_debugaccess;
  wire             std_2s60_burst_7_upstream_read;
  wire    [ 31: 0] std_2s60_burst_7_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_7_upstream_readdata_from_sa;
  wire             std_2s60_burst_7_upstream_readdatavalid;
  wire             std_2s60_burst_7_upstream_waitrequest;
  wire             std_2s60_burst_7_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_7_upstream_write;
  wire    [ 31: 0] std_2s60_burst_7_upstream_writedata;
  wire    [ 15: 0] std_2s60_burst_8_downstream_address;
  wire    [ 15: 0] std_2s60_burst_8_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_8_downstream_arbitrationshare;
  wire             std_2s60_burst_8_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_8_downstream_byteenable;
  wire             std_2s60_burst_8_downstream_debugaccess;
  wire             std_2s60_burst_8_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_granted_lan91c111_s1;
  wire    [  1: 0] std_2s60_burst_8_downstream_latency_counter;
  wire    [ 15: 0] std_2s60_burst_8_downstream_nativeaddress;
  wire             std_2s60_burst_8_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_read;
  wire             std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1;
  wire    [ 31: 0] std_2s60_burst_8_downstream_readdata;
  wire             std_2s60_burst_8_downstream_readdatavalid;
  wire             std_2s60_burst_8_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_8_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_8_downstream_reset_n;
  wire             std_2s60_burst_8_downstream_waitrequest;
  wire             std_2s60_burst_8_downstream_write;
  wire    [ 31: 0] std_2s60_burst_8_downstream_writedata;
  wire    [ 15: 0] std_2s60_burst_8_upstream_address;
  wire    [ 17: 0] std_2s60_burst_8_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_8_upstream_byteenable;
  wire             std_2s60_burst_8_upstream_debugaccess;
  wire             std_2s60_burst_8_upstream_read;
  wire    [ 31: 0] std_2s60_burst_8_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_8_upstream_readdata_from_sa;
  wire             std_2s60_burst_8_upstream_readdatavalid;
  wire             std_2s60_burst_8_upstream_waitrequest;
  wire             std_2s60_burst_8_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_8_upstream_write;
  wire    [ 31: 0] std_2s60_burst_8_upstream_writedata;
  wire    [ 15: 0] std_2s60_burst_9_downstream_address;
  wire    [ 15: 0] std_2s60_burst_9_downstream_address_to_slave;
  wire    [  3: 0] std_2s60_burst_9_downstream_arbitrationshare;
  wire             std_2s60_burst_9_downstream_burstcount;
  wire    [  3: 0] std_2s60_burst_9_downstream_byteenable;
  wire             std_2s60_burst_9_downstream_debugaccess;
  wire             std_2s60_burst_9_downstream_granted_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_granted_lan91c111_s1;
  wire    [  1: 0] std_2s60_burst_9_downstream_latency_counter;
  wire    [ 15: 0] std_2s60_burst_9_downstream_nativeaddress;
  wire             std_2s60_burst_9_downstream_qualified_request_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_qualified_request_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_read;
  wire             std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1;
  wire    [ 31: 0] std_2s60_burst_9_downstream_readdata;
  wire             std_2s60_burst_9_downstream_readdatavalid;
  wire             std_2s60_burst_9_downstream_requests_ext_ram_s1;
  wire             std_2s60_burst_9_downstream_requests_lan91c111_s1;
  wire             std_2s60_burst_9_downstream_reset_n;
  wire             std_2s60_burst_9_downstream_waitrequest;
  wire             std_2s60_burst_9_downstream_write;
  wire    [ 31: 0] std_2s60_burst_9_downstream_writedata;
  wire    [ 15: 0] std_2s60_burst_9_upstream_address;
  wire    [  3: 0] std_2s60_burst_9_upstream_burstcount;
  wire    [ 17: 0] std_2s60_burst_9_upstream_byteaddress;
  wire    [  3: 0] std_2s60_burst_9_upstream_byteenable;
  wire             std_2s60_burst_9_upstream_debugaccess;
  wire             std_2s60_burst_9_upstream_read;
  wire    [ 31: 0] std_2s60_burst_9_upstream_readdata;
  wire    [ 31: 0] std_2s60_burst_9_upstream_readdata_from_sa;
  wire             std_2s60_burst_9_upstream_readdatavalid;
  wire             std_2s60_burst_9_upstream_waitrequest;
  wire             std_2s60_burst_9_upstream_waitrequest_from_sa;
  wire             std_2s60_burst_9_upstream_write;
  wire    [ 31: 0] std_2s60_burst_9_upstream_writedata;
  wire    [  2: 0] sys_clk_timer_s1_address;
  wire             sys_clk_timer_s1_chipselect;
  wire             sys_clk_timer_s1_irq;
  wire             sys_clk_timer_s1_irq_from_sa;
  wire    [ 15: 0] sys_clk_timer_s1_readdata;
  wire    [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  wire             sys_clk_timer_s1_reset_n;
  wire             sys_clk_timer_s1_write_n;
  wire    [ 15: 0] sys_clk_timer_s1_writedata;
  wire             sysid_control_slave_address;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             write_n_to_the_ext_flash;
  wire             write_n_to_the_ext_ram;
  wire    [ 11: 0] zs_addr_from_the_sdram;
  wire    [  1: 0] zs_ba_from_the_sdram;
  wire             zs_cas_n_from_the_sdram;
  wire             zs_cke_from_the_sdram;
  wire             zs_cs_n_from_the_sdram;
  wire    [ 31: 0] zs_dq_to_and_from_the_sdram;
  wire    [  3: 0] zs_dqm_from_the_sdram;
  wire             zs_ras_n_from_the_sdram;
  wire             zs_we_n_from_the_sdram;
  ad_buf_s1_arbitrator the_ad_buf_s1
    (
      .ad_buf_s1_address                                        (ad_buf_s1_address),
      .ad_buf_s1_chipselect_n                                   (ad_buf_s1_chipselect_n),
      .ad_buf_s1_read                                           (ad_buf_s1_read),
      .ad_buf_s1_readdata                                       (ad_buf_s1_readdata),
      .ad_buf_s1_readdata_from_sa                               (ad_buf_s1_readdata_from_sa),
      .ad_buf_s1_reset_n                                        (ad_buf_s1_reset_n),
      .ad_buf_s1_waitrequest                                    (ad_buf_s1_waitrequest),
      .ad_buf_s1_waitrequest_from_sa                            (ad_buf_s1_waitrequest_from_sa),
      .clk                                                      (clk),
      .d1_ad_buf_s1_end_xfer                                    (d1_ad_buf_s1_end_xfer),
      .reset_n                                                  (clk_reset_n),
      .std_2s60_burst_17_downstream_address_to_slave            (std_2s60_burst_17_downstream_address_to_slave),
      .std_2s60_burst_17_downstream_arbitrationshare            (std_2s60_burst_17_downstream_arbitrationshare),
      .std_2s60_burst_17_downstream_burstcount                  (std_2s60_burst_17_downstream_burstcount),
      .std_2s60_burst_17_downstream_granted_ad_buf_s1           (std_2s60_burst_17_downstream_granted_ad_buf_s1),
      .std_2s60_burst_17_downstream_latency_counter             (std_2s60_burst_17_downstream_latency_counter),
      .std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 (std_2s60_burst_17_downstream_qualified_request_ad_buf_s1),
      .std_2s60_burst_17_downstream_read                        (std_2s60_burst_17_downstream_read),
      .std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1   (std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1),
      .std_2s60_burst_17_downstream_requests_ad_buf_s1          (std_2s60_burst_17_downstream_requests_ad_buf_s1),
      .std_2s60_burst_17_downstream_write                       (std_2s60_burst_17_downstream_write),
      .std_2s60_burst_18_downstream_address_to_slave            (std_2s60_burst_18_downstream_address_to_slave),
      .std_2s60_burst_18_downstream_arbitrationshare            (std_2s60_burst_18_downstream_arbitrationshare),
      .std_2s60_burst_18_downstream_burstcount                  (std_2s60_burst_18_downstream_burstcount),
      .std_2s60_burst_18_downstream_granted_ad_buf_s1           (std_2s60_burst_18_downstream_granted_ad_buf_s1),
      .std_2s60_burst_18_downstream_latency_counter             (std_2s60_burst_18_downstream_latency_counter),
      .std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 (std_2s60_burst_18_downstream_qualified_request_ad_buf_s1),
      .std_2s60_burst_18_downstream_read                        (std_2s60_burst_18_downstream_read),
      .std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1   (std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1),
      .std_2s60_burst_18_downstream_requests_ad_buf_s1          (std_2s60_burst_18_downstream_requests_ad_buf_s1),
      .std_2s60_burst_18_downstream_write                       (std_2s60_burst_18_downstream_write)
    );

  ad_buf the_ad_buf
    (
      .a2dc    (a2dc_to_the_ad_buf),
      .a2do    (ad_buf_s1_readdata),
      .adclk   (adclk_to_the_ad_buf),
      .addr    (ad_buf_s1_address),
      .cs_n    (ad_buf_s1_chipselect_n),
      .rd      (ad_buf_s1_read),
      .rdclk   (clk),
      .rst_n   (ad_buf_s1_reset_n),
      .waitreq (ad_buf_s1_waitrequest),
      .wrclk   (wrclk_to_the_ad_buf)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                                 (clk),
      .cpu_jtag_debug_module_address                                       (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                                 (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                                    (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                                    (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                                   (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                      (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                              (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset                                         (cpu_jtag_debug_module_reset),
      .cpu_jtag_debug_module_reset_n                                       (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                                  (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                          (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                         (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                     (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                                   (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                             (clk_reset_n),
      .std_2s60_burst_0_downstream_address_to_slave                        (std_2s60_burst_0_downstream_address_to_slave),
      .std_2s60_burst_0_downstream_arbitrationshare                        (std_2s60_burst_0_downstream_arbitrationshare),
      .std_2s60_burst_0_downstream_burstcount                              (std_2s60_burst_0_downstream_burstcount),
      .std_2s60_burst_0_downstream_byteenable                              (std_2s60_burst_0_downstream_byteenable),
      .std_2s60_burst_0_downstream_debugaccess                             (std_2s60_burst_0_downstream_debugaccess),
      .std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module           (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_latency_counter                         (std_2s60_burst_0_downstream_latency_counter),
      .std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module (std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_read                                    (std_2s60_burst_0_downstream_read),
      .std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module   (std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module          (std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_write                                   (std_2s60_burst_0_downstream_write),
      .std_2s60_burst_0_downstream_writedata                               (std_2s60_burst_0_downstream_writedata),
      .std_2s60_burst_1_downstream_address_to_slave                        (std_2s60_burst_1_downstream_address_to_slave),
      .std_2s60_burst_1_downstream_arbitrationshare                        (std_2s60_burst_1_downstream_arbitrationshare),
      .std_2s60_burst_1_downstream_burstcount                              (std_2s60_burst_1_downstream_burstcount),
      .std_2s60_burst_1_downstream_byteenable                              (std_2s60_burst_1_downstream_byteenable),
      .std_2s60_burst_1_downstream_debugaccess                             (std_2s60_burst_1_downstream_debugaccess),
      .std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module           (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_latency_counter                         (std_2s60_burst_1_downstream_latency_counter),
      .std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module (std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_read                                    (std_2s60_burst_1_downstream_read),
      .std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module   (std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module          (std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_write                                   (std_2s60_burst_1_downstream_write),
      .std_2s60_burst_1_downstream_writedata                               (std_2s60_burst_1_downstream_writedata)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .clk                                                                       (clk),
      .cpu_data_master_address                                                   (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_byteenable_std_2s60_burst_3_upstream                      (cpu_data_master_byteenable_std_2s60_burst_3_upstream),
      .cpu_data_master_dbs_address                                               (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_8                                               (cpu_data_master_dbs_write_8),
      .cpu_data_master_granted_std_2s60_burst_10_upstream                        (cpu_data_master_granted_std_2s60_burst_10_upstream),
      .cpu_data_master_granted_std_2s60_burst_11_upstream                        (cpu_data_master_granted_std_2s60_burst_11_upstream),
      .cpu_data_master_granted_std_2s60_burst_12_upstream                        (cpu_data_master_granted_std_2s60_burst_12_upstream),
      .cpu_data_master_granted_std_2s60_burst_13_upstream                        (cpu_data_master_granted_std_2s60_burst_13_upstream),
      .cpu_data_master_granted_std_2s60_burst_14_upstream                        (cpu_data_master_granted_std_2s60_burst_14_upstream),
      .cpu_data_master_granted_std_2s60_burst_16_upstream                        (cpu_data_master_granted_std_2s60_burst_16_upstream),
      .cpu_data_master_granted_std_2s60_burst_17_upstream                        (cpu_data_master_granted_std_2s60_burst_17_upstream),
      .cpu_data_master_granted_std_2s60_burst_1_upstream                         (cpu_data_master_granted_std_2s60_burst_1_upstream),
      .cpu_data_master_granted_std_2s60_burst_3_upstream                         (cpu_data_master_granted_std_2s60_burst_3_upstream),
      .cpu_data_master_granted_std_2s60_burst_5_upstream                         (cpu_data_master_granted_std_2s60_burst_5_upstream),
      .cpu_data_master_granted_std_2s60_burst_7_upstream                         (cpu_data_master_granted_std_2s60_burst_7_upstream),
      .cpu_data_master_granted_std_2s60_burst_9_upstream                         (cpu_data_master_granted_std_2s60_burst_9_upstream),
      .cpu_data_master_irq                                                       (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_10_upstream              (cpu_data_master_qualified_request_std_2s60_burst_10_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_11_upstream              (cpu_data_master_qualified_request_std_2s60_burst_11_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_12_upstream              (cpu_data_master_qualified_request_std_2s60_burst_12_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_13_upstream              (cpu_data_master_qualified_request_std_2s60_burst_13_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_14_upstream              (cpu_data_master_qualified_request_std_2s60_burst_14_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_16_upstream              (cpu_data_master_qualified_request_std_2s60_burst_16_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_17_upstream              (cpu_data_master_qualified_request_std_2s60_burst_17_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_1_upstream               (cpu_data_master_qualified_request_std_2s60_burst_1_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_3_upstream               (cpu_data_master_qualified_request_std_2s60_burst_3_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_5_upstream               (cpu_data_master_qualified_request_std_2s60_burst_5_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_7_upstream               (cpu_data_master_qualified_request_std_2s60_burst_7_upstream),
      .cpu_data_master_qualified_request_std_2s60_burst_9_upstream               (cpu_data_master_qualified_request_std_2s60_burst_9_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_readdata                                                  (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                             (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_std_2s60_burst_10_upstream                       (cpu_data_master_requests_std_2s60_burst_10_upstream),
      .cpu_data_master_requests_std_2s60_burst_11_upstream                       (cpu_data_master_requests_std_2s60_burst_11_upstream),
      .cpu_data_master_requests_std_2s60_burst_12_upstream                       (cpu_data_master_requests_std_2s60_burst_12_upstream),
      .cpu_data_master_requests_std_2s60_burst_13_upstream                       (cpu_data_master_requests_std_2s60_burst_13_upstream),
      .cpu_data_master_requests_std_2s60_burst_14_upstream                       (cpu_data_master_requests_std_2s60_burst_14_upstream),
      .cpu_data_master_requests_std_2s60_burst_16_upstream                       (cpu_data_master_requests_std_2s60_burst_16_upstream),
      .cpu_data_master_requests_std_2s60_burst_17_upstream                       (cpu_data_master_requests_std_2s60_burst_17_upstream),
      .cpu_data_master_requests_std_2s60_burst_1_upstream                        (cpu_data_master_requests_std_2s60_burst_1_upstream),
      .cpu_data_master_requests_std_2s60_burst_3_upstream                        (cpu_data_master_requests_std_2s60_burst_3_upstream),
      .cpu_data_master_requests_std_2s60_burst_5_upstream                        (cpu_data_master_requests_std_2s60_burst_5_upstream),
      .cpu_data_master_requests_std_2s60_burst_7_upstream                        (cpu_data_master_requests_std_2s60_burst_7_upstream),
      .cpu_data_master_requests_std_2s60_burst_9_upstream                        (cpu_data_master_requests_std_2s60_burst_9_upstream),
      .cpu_data_master_waitrequest                                               (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_irq_from_the_lan91c111                                                 (d1_irq_from_the_lan91c111),
      .d1_std_2s60_burst_10_upstream_end_xfer                                    (d1_std_2s60_burst_10_upstream_end_xfer),
      .d1_std_2s60_burst_11_upstream_end_xfer                                    (d1_std_2s60_burst_11_upstream_end_xfer),
      .d1_std_2s60_burst_12_upstream_end_xfer                                    (d1_std_2s60_burst_12_upstream_end_xfer),
      .d1_std_2s60_burst_13_upstream_end_xfer                                    (d1_std_2s60_burst_13_upstream_end_xfer),
      .d1_std_2s60_burst_14_upstream_end_xfer                                    (d1_std_2s60_burst_14_upstream_end_xfer),
      .d1_std_2s60_burst_16_upstream_end_xfer                                    (d1_std_2s60_burst_16_upstream_end_xfer),
      .d1_std_2s60_burst_17_upstream_end_xfer                                    (d1_std_2s60_burst_17_upstream_end_xfer),
      .d1_std_2s60_burst_1_upstream_end_xfer                                     (d1_std_2s60_burst_1_upstream_end_xfer),
      .d1_std_2s60_burst_3_upstream_end_xfer                                     (d1_std_2s60_burst_3_upstream_end_xfer),
      .d1_std_2s60_burst_5_upstream_end_xfer                                     (d1_std_2s60_burst_5_upstream_end_xfer),
      .d1_std_2s60_burst_7_upstream_end_xfer                                     (d1_std_2s60_burst_7_upstream_end_xfer),
      .d1_std_2s60_burst_9_upstream_end_xfer                                     (d1_std_2s60_burst_9_upstream_end_xfer),
      .high_res_timer_s1_irq_from_sa                                             (high_res_timer_s1_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                   (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_10_upstream_readdata_from_sa                               (std_2s60_burst_10_upstream_readdata_from_sa),
      .std_2s60_burst_10_upstream_waitrequest_from_sa                            (std_2s60_burst_10_upstream_waitrequest_from_sa),
      .std_2s60_burst_11_upstream_readdata_from_sa                               (std_2s60_burst_11_upstream_readdata_from_sa),
      .std_2s60_burst_11_upstream_waitrequest_from_sa                            (std_2s60_burst_11_upstream_waitrequest_from_sa),
      .std_2s60_burst_12_upstream_readdata_from_sa                               (std_2s60_burst_12_upstream_readdata_from_sa),
      .std_2s60_burst_12_upstream_waitrequest_from_sa                            (std_2s60_burst_12_upstream_waitrequest_from_sa),
      .std_2s60_burst_13_upstream_readdata_from_sa                               (std_2s60_burst_13_upstream_readdata_from_sa),
      .std_2s60_burst_13_upstream_waitrequest_from_sa                            (std_2s60_burst_13_upstream_waitrequest_from_sa),
      .std_2s60_burst_14_upstream_readdata_from_sa                               (std_2s60_burst_14_upstream_readdata_from_sa),
      .std_2s60_burst_14_upstream_waitrequest_from_sa                            (std_2s60_burst_14_upstream_waitrequest_from_sa),
      .std_2s60_burst_16_upstream_readdata_from_sa                               (std_2s60_burst_16_upstream_readdata_from_sa),
      .std_2s60_burst_16_upstream_waitrequest_from_sa                            (std_2s60_burst_16_upstream_waitrequest_from_sa),
      .std_2s60_burst_17_upstream_readdata_from_sa                               (std_2s60_burst_17_upstream_readdata_from_sa),
      .std_2s60_burst_17_upstream_waitrequest_from_sa                            (std_2s60_burst_17_upstream_waitrequest_from_sa),
      .std_2s60_burst_1_upstream_readdata_from_sa                                (std_2s60_burst_1_upstream_readdata_from_sa),
      .std_2s60_burst_1_upstream_waitrequest_from_sa                             (std_2s60_burst_1_upstream_waitrequest_from_sa),
      .std_2s60_burst_3_upstream_readdata_from_sa                                (std_2s60_burst_3_upstream_readdata_from_sa),
      .std_2s60_burst_3_upstream_waitrequest_from_sa                             (std_2s60_burst_3_upstream_waitrequest_from_sa),
      .std_2s60_burst_5_upstream_readdata_from_sa                                (std_2s60_burst_5_upstream_readdata_from_sa),
      .std_2s60_burst_5_upstream_waitrequest_from_sa                             (std_2s60_burst_5_upstream_waitrequest_from_sa),
      .std_2s60_burst_7_upstream_readdata_from_sa                                (std_2s60_burst_7_upstream_readdata_from_sa),
      .std_2s60_burst_7_upstream_waitrequest_from_sa                             (std_2s60_burst_7_upstream_waitrequest_from_sa),
      .std_2s60_burst_9_upstream_readdata_from_sa                                (std_2s60_burst_9_upstream_readdata_from_sa),
      .std_2s60_burst_9_upstream_waitrequest_from_sa                             (std_2s60_burst_9_upstream_waitrequest_from_sa),
      .sys_clk_timer_s1_irq_from_sa                                              (sys_clk_timer_s1_irq_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address                                                   (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_dbs_address                                               (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_std_2s60_burst_0_upstream                         (cpu_instruction_master_granted_std_2s60_burst_0_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_15_upstream                        (cpu_instruction_master_granted_std_2s60_burst_15_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_18_upstream                        (cpu_instruction_master_granted_std_2s60_burst_18_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_2_upstream                         (cpu_instruction_master_granted_std_2s60_burst_2_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_4_upstream                         (cpu_instruction_master_granted_std_2s60_burst_4_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_6_upstream                         (cpu_instruction_master_granted_std_2s60_burst_6_upstream),
      .cpu_instruction_master_granted_std_2s60_burst_8_upstream                         (cpu_instruction_master_granted_std_2s60_burst_8_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream              (cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream              (cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream),
      .cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream                (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream                (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_readdata                                                  (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                                             (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_std_2s60_burst_0_upstream                        (cpu_instruction_master_requests_std_2s60_burst_0_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_15_upstream                       (cpu_instruction_master_requests_std_2s60_burst_15_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_18_upstream                       (cpu_instruction_master_requests_std_2s60_burst_18_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_2_upstream                        (cpu_instruction_master_requests_std_2s60_burst_2_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_4_upstream                        (cpu_instruction_master_requests_std_2s60_burst_4_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_6_upstream                        (cpu_instruction_master_requests_std_2s60_burst_6_upstream),
      .cpu_instruction_master_requests_std_2s60_burst_8_upstream                        (cpu_instruction_master_requests_std_2s60_burst_8_upstream),
      .cpu_instruction_master_waitrequest                                               (cpu_instruction_master_waitrequest),
      .d1_std_2s60_burst_0_upstream_end_xfer                                            (d1_std_2s60_burst_0_upstream_end_xfer),
      .d1_std_2s60_burst_15_upstream_end_xfer                                           (d1_std_2s60_burst_15_upstream_end_xfer),
      .d1_std_2s60_burst_18_upstream_end_xfer                                           (d1_std_2s60_burst_18_upstream_end_xfer),
      .d1_std_2s60_burst_2_upstream_end_xfer                                            (d1_std_2s60_burst_2_upstream_end_xfer),
      .d1_std_2s60_burst_4_upstream_end_xfer                                            (d1_std_2s60_burst_4_upstream_end_xfer),
      .d1_std_2s60_burst_6_upstream_end_xfer                                            (d1_std_2s60_burst_6_upstream_end_xfer),
      .d1_std_2s60_burst_8_upstream_end_xfer                                            (d1_std_2s60_burst_8_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_0_upstream_readdata_from_sa                                       (std_2s60_burst_0_upstream_readdata_from_sa),
      .std_2s60_burst_0_upstream_waitrequest_from_sa                                    (std_2s60_burst_0_upstream_waitrequest_from_sa),
      .std_2s60_burst_15_upstream_readdata_from_sa                                      (std_2s60_burst_15_upstream_readdata_from_sa),
      .std_2s60_burst_15_upstream_waitrequest_from_sa                                   (std_2s60_burst_15_upstream_waitrequest_from_sa),
      .std_2s60_burst_18_upstream_readdata_from_sa                                      (std_2s60_burst_18_upstream_readdata_from_sa),
      .std_2s60_burst_18_upstream_waitrequest_from_sa                                   (std_2s60_burst_18_upstream_waitrequest_from_sa),
      .std_2s60_burst_2_upstream_readdata_from_sa                                       (std_2s60_burst_2_upstream_readdata_from_sa),
      .std_2s60_burst_2_upstream_waitrequest_from_sa                                    (std_2s60_burst_2_upstream_waitrequest_from_sa),
      .std_2s60_burst_4_upstream_readdata_from_sa                                       (std_2s60_burst_4_upstream_readdata_from_sa),
      .std_2s60_burst_4_upstream_waitrequest_from_sa                                    (std_2s60_burst_4_upstream_waitrequest_from_sa),
      .std_2s60_burst_6_upstream_readdata_from_sa                                       (std_2s60_burst_6_upstream_readdata_from_sa),
      .std_2s60_burst_6_upstream_waitrequest_from_sa                                    (std_2s60_burst_6_upstream_waitrequest_from_sa),
      .std_2s60_burst_8_upstream_readdata_from_sa                                       (std_2s60_burst_8_upstream_readdata_from_sa),
      .std_2s60_burst_8_upstream_waitrequest_from_sa                                    (std_2s60_burst_8_upstream_waitrequest_from_sa)
    );

  cpu the_cpu
    (
      .clk                                   (clk),
      .d_address                             (cpu_data_master_address),
      .d_burstcount                          (cpu_data_master_burstcount),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_burstcount                          (cpu_instruction_master_burstcount),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_clk                 (clk),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_reset               (cpu_jtag_debug_module_reset),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  ext_flash_bus_avalon_slave_arbitrator the_ext_flash_bus_avalon_slave
    (
      .clk                                                        (clk),
      .d1_ext_flash_bus_avalon_slave_end_xfer                     (d1_ext_flash_bus_avalon_slave_end_xfer),
      .ext_flash_bus_address                                      (ext_flash_bus_address),
      .ext_flash_bus_data                                         (ext_flash_bus_data),
      .ext_flash_bus_readn                                        (ext_flash_bus_readn),
      .ext_flash_s1_wait_counter_eq_0                             (ext_flash_s1_wait_counter_eq_0),
      .incoming_ext_flash_bus_data_with_Xs_converted_to_0         (incoming_ext_flash_bus_data_with_Xs_converted_to_0),
      .reset_n                                                    (clk_reset_n),
      .select_n_to_the_ext_flash                                  (select_n_to_the_ext_flash),
      .std_2s60_burst_2_downstream_address_to_slave               (std_2s60_burst_2_downstream_address_to_slave),
      .std_2s60_burst_2_downstream_arbitrationshare               (std_2s60_burst_2_downstream_arbitrationshare),
      .std_2s60_burst_2_downstream_burstcount                     (std_2s60_burst_2_downstream_burstcount),
      .std_2s60_burst_2_downstream_byteenable                     (std_2s60_burst_2_downstream_byteenable),
      .std_2s60_burst_2_downstream_granted_ext_flash_s1           (std_2s60_burst_2_downstream_granted_ext_flash_s1),
      .std_2s60_burst_2_downstream_latency_counter                (std_2s60_burst_2_downstream_latency_counter),
      .std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 (std_2s60_burst_2_downstream_qualified_request_ext_flash_s1),
      .std_2s60_burst_2_downstream_read                           (std_2s60_burst_2_downstream_read),
      .std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1   (std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1),
      .std_2s60_burst_2_downstream_requests_ext_flash_s1          (std_2s60_burst_2_downstream_requests_ext_flash_s1),
      .std_2s60_burst_2_downstream_write                          (std_2s60_burst_2_downstream_write),
      .std_2s60_burst_2_downstream_writedata                      (std_2s60_burst_2_downstream_writedata),
      .std_2s60_burst_3_downstream_address_to_slave               (std_2s60_burst_3_downstream_address_to_slave),
      .std_2s60_burst_3_downstream_arbitrationshare               (std_2s60_burst_3_downstream_arbitrationshare),
      .std_2s60_burst_3_downstream_burstcount                     (std_2s60_burst_3_downstream_burstcount),
      .std_2s60_burst_3_downstream_byteenable                     (std_2s60_burst_3_downstream_byteenable),
      .std_2s60_burst_3_downstream_granted_ext_flash_s1           (std_2s60_burst_3_downstream_granted_ext_flash_s1),
      .std_2s60_burst_3_downstream_latency_counter                (std_2s60_burst_3_downstream_latency_counter),
      .std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 (std_2s60_burst_3_downstream_qualified_request_ext_flash_s1),
      .std_2s60_burst_3_downstream_read                           (std_2s60_burst_3_downstream_read),
      .std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1   (std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1),
      .std_2s60_burst_3_downstream_requests_ext_flash_s1          (std_2s60_burst_3_downstream_requests_ext_flash_s1),
      .std_2s60_burst_3_downstream_write                          (std_2s60_burst_3_downstream_write),
      .std_2s60_burst_3_downstream_writedata                      (std_2s60_burst_3_downstream_writedata),
      .write_n_to_the_ext_flash                                   (write_n_to_the_ext_flash)
    );

  ext_ram_bus_avalon_slave_arbitrator the_ext_ram_bus_avalon_slave
    (
      .be_n_to_the_ext_ram                                        (be_n_to_the_ext_ram),
      .clk                                                        (clk),
      .d1_ext_ram_bus_avalon_slave_end_xfer                       (d1_ext_ram_bus_avalon_slave_end_xfer),
      .d1_irq_from_the_lan91c111                                  (d1_irq_from_the_lan91c111),
      .ext_ram_bus_address                                        (ext_ram_bus_address),
      .ext_ram_bus_byteenablen                                    (ext_ram_bus_byteenablen),
      .ext_ram_bus_data                                           (ext_ram_bus_data),
      .ext_ram_s1_wait_counter_eq_0                               (ext_ram_s1_wait_counter_eq_0),
      .incoming_ext_ram_bus_data                                  (incoming_ext_ram_bus_data),
      .ior_n_to_the_lan91c111                                     (ior_n_to_the_lan91c111),
      .iow_n_to_the_lan91c111                                     (iow_n_to_the_lan91c111),
      .irq_from_the_lan91c111                                     (irq_from_the_lan91c111),
      .lan91c111_s1_wait_counter_eq_0                             (lan91c111_s1_wait_counter_eq_0),
      .read_n_to_the_ext_ram                                      (read_n_to_the_ext_ram),
      .reset_n                                                    (clk_reset_n),
      .reset_to_the_lan91c111                                     (reset_to_the_lan91c111),
      .select_n_to_the_ext_ram                                    (select_n_to_the_ext_ram),
      .std_2s60_burst_4_downstream_address_to_slave               (std_2s60_burst_4_downstream_address_to_slave),
      .std_2s60_burst_4_downstream_arbitrationshare               (std_2s60_burst_4_downstream_arbitrationshare),
      .std_2s60_burst_4_downstream_burstcount                     (std_2s60_burst_4_downstream_burstcount),
      .std_2s60_burst_4_downstream_byteenable                     (std_2s60_burst_4_downstream_byteenable),
      .std_2s60_burst_4_downstream_granted_ext_ram_s1             (std_2s60_burst_4_downstream_granted_ext_ram_s1),
      .std_2s60_burst_4_downstream_granted_lan91c111_s1           (std_2s60_burst_4_downstream_granted_lan91c111_s1),
      .std_2s60_burst_4_downstream_latency_counter                (std_2s60_burst_4_downstream_latency_counter),
      .std_2s60_burst_4_downstream_nativeaddress                  (std_2s60_burst_4_downstream_nativeaddress),
      .std_2s60_burst_4_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_4_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_4_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_4_downstream_read                           (std_2s60_burst_4_downstream_read),
      .std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_4_downstream_requests_ext_ram_s1            (std_2s60_burst_4_downstream_requests_ext_ram_s1),
      .std_2s60_burst_4_downstream_requests_lan91c111_s1          (std_2s60_burst_4_downstream_requests_lan91c111_s1),
      .std_2s60_burst_4_downstream_write                          (std_2s60_burst_4_downstream_write),
      .std_2s60_burst_4_downstream_writedata                      (std_2s60_burst_4_downstream_writedata),
      .std_2s60_burst_5_downstream_address_to_slave               (std_2s60_burst_5_downstream_address_to_slave),
      .std_2s60_burst_5_downstream_arbitrationshare               (std_2s60_burst_5_downstream_arbitrationshare),
      .std_2s60_burst_5_downstream_burstcount                     (std_2s60_burst_5_downstream_burstcount),
      .std_2s60_burst_5_downstream_byteenable                     (std_2s60_burst_5_downstream_byteenable),
      .std_2s60_burst_5_downstream_granted_ext_ram_s1             (std_2s60_burst_5_downstream_granted_ext_ram_s1),
      .std_2s60_burst_5_downstream_granted_lan91c111_s1           (std_2s60_burst_5_downstream_granted_lan91c111_s1),
      .std_2s60_burst_5_downstream_latency_counter                (std_2s60_burst_5_downstream_latency_counter),
      .std_2s60_burst_5_downstream_nativeaddress                  (std_2s60_burst_5_downstream_nativeaddress),
      .std_2s60_burst_5_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_5_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_5_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_5_downstream_read                           (std_2s60_burst_5_downstream_read),
      .std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_5_downstream_requests_ext_ram_s1            (std_2s60_burst_5_downstream_requests_ext_ram_s1),
      .std_2s60_burst_5_downstream_requests_lan91c111_s1          (std_2s60_burst_5_downstream_requests_lan91c111_s1),
      .std_2s60_burst_5_downstream_write                          (std_2s60_burst_5_downstream_write),
      .std_2s60_burst_5_downstream_writedata                      (std_2s60_burst_5_downstream_writedata),
      .std_2s60_burst_8_downstream_address_to_slave               (std_2s60_burst_8_downstream_address_to_slave),
      .std_2s60_burst_8_downstream_arbitrationshare               (std_2s60_burst_8_downstream_arbitrationshare),
      .std_2s60_burst_8_downstream_burstcount                     (std_2s60_burst_8_downstream_burstcount),
      .std_2s60_burst_8_downstream_byteenable                     (std_2s60_burst_8_downstream_byteenable),
      .std_2s60_burst_8_downstream_granted_ext_ram_s1             (std_2s60_burst_8_downstream_granted_ext_ram_s1),
      .std_2s60_burst_8_downstream_granted_lan91c111_s1           (std_2s60_burst_8_downstream_granted_lan91c111_s1),
      .std_2s60_burst_8_downstream_latency_counter                (std_2s60_burst_8_downstream_latency_counter),
      .std_2s60_burst_8_downstream_nativeaddress                  (std_2s60_burst_8_downstream_nativeaddress),
      .std_2s60_burst_8_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_8_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_8_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_8_downstream_read                           (std_2s60_burst_8_downstream_read),
      .std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_8_downstream_requests_ext_ram_s1            (std_2s60_burst_8_downstream_requests_ext_ram_s1),
      .std_2s60_burst_8_downstream_requests_lan91c111_s1          (std_2s60_burst_8_downstream_requests_lan91c111_s1),
      .std_2s60_burst_8_downstream_write                          (std_2s60_burst_8_downstream_write),
      .std_2s60_burst_8_downstream_writedata                      (std_2s60_burst_8_downstream_writedata),
      .std_2s60_burst_9_downstream_address_to_slave               (std_2s60_burst_9_downstream_address_to_slave),
      .std_2s60_burst_9_downstream_arbitrationshare               (std_2s60_burst_9_downstream_arbitrationshare),
      .std_2s60_burst_9_downstream_burstcount                     (std_2s60_burst_9_downstream_burstcount),
      .std_2s60_burst_9_downstream_byteenable                     (std_2s60_burst_9_downstream_byteenable),
      .std_2s60_burst_9_downstream_granted_ext_ram_s1             (std_2s60_burst_9_downstream_granted_ext_ram_s1),
      .std_2s60_burst_9_downstream_granted_lan91c111_s1           (std_2s60_burst_9_downstream_granted_lan91c111_s1),
      .std_2s60_burst_9_downstream_latency_counter                (std_2s60_burst_9_downstream_latency_counter),
      .std_2s60_burst_9_downstream_nativeaddress                  (std_2s60_burst_9_downstream_nativeaddress),
      .std_2s60_burst_9_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_9_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_9_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_9_downstream_read                           (std_2s60_burst_9_downstream_read),
      .std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_9_downstream_requests_ext_ram_s1            (std_2s60_burst_9_downstream_requests_ext_ram_s1),
      .std_2s60_burst_9_downstream_requests_lan91c111_s1          (std_2s60_burst_9_downstream_requests_lan91c111_s1),
      .std_2s60_burst_9_downstream_write                          (std_2s60_burst_9_downstream_write),
      .std_2s60_burst_9_downstream_writedata                      (std_2s60_burst_9_downstream_writedata),
      .write_n_to_the_ext_ram                                     (write_n_to_the_ext_ram)
    );

  high_res_timer_s1_arbitrator the_high_res_timer_s1
    (
      .clk                                                              (clk),
      .d1_high_res_timer_s1_end_xfer                                    (d1_high_res_timer_s1_end_xfer),
      .high_res_timer_s1_address                                        (high_res_timer_s1_address),
      .high_res_timer_s1_chipselect                                     (high_res_timer_s1_chipselect),
      .high_res_timer_s1_irq                                            (high_res_timer_s1_irq),
      .high_res_timer_s1_irq_from_sa                                    (high_res_timer_s1_irq_from_sa),
      .high_res_timer_s1_readdata                                       (high_res_timer_s1_readdata),
      .high_res_timer_s1_readdata_from_sa                               (high_res_timer_s1_readdata_from_sa),
      .high_res_timer_s1_reset_n                                        (high_res_timer_s1_reset_n),
      .high_res_timer_s1_write_n                                        (high_res_timer_s1_write_n),
      .high_res_timer_s1_writedata                                      (high_res_timer_s1_writedata),
      .reset_n                                                          (clk_reset_n),
      .std_2s60_burst_12_downstream_address_to_slave                    (std_2s60_burst_12_downstream_address_to_slave),
      .std_2s60_burst_12_downstream_arbitrationshare                    (std_2s60_burst_12_downstream_arbitrationshare),
      .std_2s60_burst_12_downstream_burstcount                          (std_2s60_burst_12_downstream_burstcount),
      .std_2s60_burst_12_downstream_granted_high_res_timer_s1           (std_2s60_burst_12_downstream_granted_high_res_timer_s1),
      .std_2s60_burst_12_downstream_latency_counter                     (std_2s60_burst_12_downstream_latency_counter),
      .std_2s60_burst_12_downstream_nativeaddress                       (std_2s60_burst_12_downstream_nativeaddress),
      .std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 (std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1),
      .std_2s60_burst_12_downstream_read                                (std_2s60_burst_12_downstream_read),
      .std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1   (std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1),
      .std_2s60_burst_12_downstream_requests_high_res_timer_s1          (std_2s60_burst_12_downstream_requests_high_res_timer_s1),
      .std_2s60_burst_12_downstream_write                               (std_2s60_burst_12_downstream_write),
      .std_2s60_burst_12_downstream_writedata                           (std_2s60_burst_12_downstream_writedata)
    );

  high_res_timer the_high_res_timer
    (
      .address    (high_res_timer_s1_address),
      .chipselect (high_res_timer_s1_chipselect),
      .clk        (clk),
      .irq        (high_res_timer_s1_irq),
      .readdata   (high_res_timer_s1_readdata),
      .reset_n    (high_res_timer_s1_reset_n),
      .write_n    (high_res_timer_s1_write_n),
      .writedata  (high_res_timer_s1_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                                        (clk),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                    (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                                        (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                                     (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                                  (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa                          (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                                            (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                    (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                                         (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                                       (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                               (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                                   (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa                           (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                                        (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                                    (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                            (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                                        (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                                      (jtag_uart_avalon_jtag_slave_writedata),
      .reset_n                                                                    (clk_reset_n),
      .std_2s60_burst_11_downstream_address_to_slave                              (std_2s60_burst_11_downstream_address_to_slave),
      .std_2s60_burst_11_downstream_arbitrationshare                              (std_2s60_burst_11_downstream_arbitrationshare),
      .std_2s60_burst_11_downstream_burstcount                                    (std_2s60_burst_11_downstream_burstcount),
      .std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave           (std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_latency_counter                               (std_2s60_burst_11_downstream_latency_counter),
      .std_2s60_burst_11_downstream_nativeaddress                                 (std_2s60_burst_11_downstream_nativeaddress),
      .std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave (std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_read                                          (std_2s60_burst_11_downstream_read),
      .std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave   (std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave          (std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_write                                         (std_2s60_burst_11_downstream_write),
      .std_2s60_burst_11_downstream_writedata                                     (std_2s60_burst_11_downstream_writedata)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (clk),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  onchip_ram_64_kbytes_s1_arbitrator the_onchip_ram_64_kbytes_s1
    (
      .clk                                                                   (clk),
      .d1_onchip_ram_64_kbytes_s1_end_xfer                                   (d1_onchip_ram_64_kbytes_s1_end_xfer),
      .onchip_ram_64_kbytes_s1_address                                       (onchip_ram_64_kbytes_s1_address),
      .onchip_ram_64_kbytes_s1_byteenable                                    (onchip_ram_64_kbytes_s1_byteenable),
      .onchip_ram_64_kbytes_s1_chipselect                                    (onchip_ram_64_kbytes_s1_chipselect),
      .onchip_ram_64_kbytes_s1_clken                                         (onchip_ram_64_kbytes_s1_clken),
      .onchip_ram_64_kbytes_s1_readdata                                      (onchip_ram_64_kbytes_s1_readdata),
      .onchip_ram_64_kbytes_s1_readdata_from_sa                              (onchip_ram_64_kbytes_s1_readdata_from_sa),
      .onchip_ram_64_kbytes_s1_write                                         (onchip_ram_64_kbytes_s1_write),
      .onchip_ram_64_kbytes_s1_writedata                                     (onchip_ram_64_kbytes_s1_writedata),
      .reset_n                                                               (clk_reset_n),
      .std_2s60_burst_6_downstream_address_to_slave                          (std_2s60_burst_6_downstream_address_to_slave),
      .std_2s60_burst_6_downstream_arbitrationshare                          (std_2s60_burst_6_downstream_arbitrationshare),
      .std_2s60_burst_6_downstream_burstcount                                (std_2s60_burst_6_downstream_burstcount),
      .std_2s60_burst_6_downstream_byteenable                                (std_2s60_burst_6_downstream_byteenable),
      .std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1           (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_latency_counter                           (std_2s60_burst_6_downstream_latency_counter),
      .std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 (std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_read                                      (std_2s60_burst_6_downstream_read),
      .std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1   (std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1          (std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_write                                     (std_2s60_burst_6_downstream_write),
      .std_2s60_burst_6_downstream_writedata                                 (std_2s60_burst_6_downstream_writedata),
      .std_2s60_burst_7_downstream_address_to_slave                          (std_2s60_burst_7_downstream_address_to_slave),
      .std_2s60_burst_7_downstream_arbitrationshare                          (std_2s60_burst_7_downstream_arbitrationshare),
      .std_2s60_burst_7_downstream_burstcount                                (std_2s60_burst_7_downstream_burstcount),
      .std_2s60_burst_7_downstream_byteenable                                (std_2s60_burst_7_downstream_byteenable),
      .std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1           (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_latency_counter                           (std_2s60_burst_7_downstream_latency_counter),
      .std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 (std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_read                                      (std_2s60_burst_7_downstream_read),
      .std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1   (std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1          (std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_write                                     (std_2s60_burst_7_downstream_write),
      .std_2s60_burst_7_downstream_writedata                                 (std_2s60_burst_7_downstream_writedata)
    );

  onchip_ram_64_kbytes the_onchip_ram_64_kbytes
    (
      .address    (onchip_ram_64_kbytes_s1_address),
      .byteenable (onchip_ram_64_kbytes_s1_byteenable),
      .chipselect (onchip_ram_64_kbytes_s1_chipselect),
      .clk        (clk),
      .clken      (onchip_ram_64_kbytes_s1_clken),
      .readdata   (onchip_ram_64_kbytes_s1_readdata),
      .write      (onchip_ram_64_kbytes_s1_write),
      .writedata  (onchip_ram_64_kbytes_s1_writedata)
    );

  reconfig_request_pio_s1_arbitrator the_reconfig_request_pio_s1
    (
      .clk                                                                    (clk),
      .d1_reconfig_request_pio_s1_end_xfer                                    (d1_reconfig_request_pio_s1_end_xfer),
      .reconfig_request_pio_s1_address                                        (reconfig_request_pio_s1_address),
      .reconfig_request_pio_s1_chipselect                                     (reconfig_request_pio_s1_chipselect),
      .reconfig_request_pio_s1_readdata                                       (reconfig_request_pio_s1_readdata),
      .reconfig_request_pio_s1_readdata_from_sa                               (reconfig_request_pio_s1_readdata_from_sa),
      .reconfig_request_pio_s1_reset_n                                        (reconfig_request_pio_s1_reset_n),
      .reconfig_request_pio_s1_write_n                                        (reconfig_request_pio_s1_write_n),
      .reconfig_request_pio_s1_writedata                                      (reconfig_request_pio_s1_writedata),
      .reset_n                                                                (clk_reset_n),
      .std_2s60_burst_13_downstream_address_to_slave                          (std_2s60_burst_13_downstream_address_to_slave),
      .std_2s60_burst_13_downstream_arbitrationshare                          (std_2s60_burst_13_downstream_arbitrationshare),
      .std_2s60_burst_13_downstream_burstcount                                (std_2s60_burst_13_downstream_burstcount),
      .std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1           (std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_latency_counter                           (std_2s60_burst_13_downstream_latency_counter),
      .std_2s60_burst_13_downstream_nativeaddress                             (std_2s60_burst_13_downstream_nativeaddress),
      .std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 (std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_read                                      (std_2s60_burst_13_downstream_read),
      .std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1   (std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1          (std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_write                                     (std_2s60_burst_13_downstream_write),
      .std_2s60_burst_13_downstream_writedata                                 (std_2s60_burst_13_downstream_writedata)
    );

  reconfig_request_pio the_reconfig_request_pio
    (
      .address    (reconfig_request_pio_s1_address),
      .bidir_port (bidir_port_to_and_from_the_reconfig_request_pio),
      .chipselect (reconfig_request_pio_s1_chipselect),
      .clk        (clk),
      .readdata   (reconfig_request_pio_s1_readdata),
      .reset_n    (reconfig_request_pio_s1_reset_n),
      .write_n    (reconfig_request_pio_s1_write_n),
      .writedata  (reconfig_request_pio_s1_writedata)
    );

  sdram_s1_arbitrator the_sdram_s1
    (
      .clk                                                                  (clk),
      .d1_sdram_s1_end_xfer                                                 (d1_sdram_s1_end_xfer),
      .reset_n                                                              (clk_reset_n),
      .sdram_s1_address                                                     (sdram_s1_address),
      .sdram_s1_byteenable_n                                                (sdram_s1_byteenable_n),
      .sdram_s1_chipselect                                                  (sdram_s1_chipselect),
      .sdram_s1_read_n                                                      (sdram_s1_read_n),
      .sdram_s1_readdata                                                    (sdram_s1_readdata),
      .sdram_s1_readdata_from_sa                                            (sdram_s1_readdata_from_sa),
      .sdram_s1_readdatavalid                                               (sdram_s1_readdatavalid),
      .sdram_s1_reset_n                                                     (sdram_s1_reset_n),
      .sdram_s1_waitrequest                                                 (sdram_s1_waitrequest),
      .sdram_s1_waitrequest_from_sa                                         (sdram_s1_waitrequest_from_sa),
      .sdram_s1_write_n                                                     (sdram_s1_write_n),
      .sdram_s1_writedata                                                   (sdram_s1_writedata),
      .std_2s60_burst_15_downstream_address_to_slave                        (std_2s60_burst_15_downstream_address_to_slave),
      .std_2s60_burst_15_downstream_arbitrationshare                        (std_2s60_burst_15_downstream_arbitrationshare),
      .std_2s60_burst_15_downstream_burstcount                              (std_2s60_burst_15_downstream_burstcount),
      .std_2s60_burst_15_downstream_byteenable                              (std_2s60_burst_15_downstream_byteenable),
      .std_2s60_burst_15_downstream_granted_sdram_s1                        (std_2s60_burst_15_downstream_granted_sdram_s1),
      .std_2s60_burst_15_downstream_latency_counter                         (std_2s60_burst_15_downstream_latency_counter),
      .std_2s60_burst_15_downstream_qualified_request_sdram_s1              (std_2s60_burst_15_downstream_qualified_request_sdram_s1),
      .std_2s60_burst_15_downstream_read                                    (std_2s60_burst_15_downstream_read),
      .std_2s60_burst_15_downstream_read_data_valid_sdram_s1                (std_2s60_burst_15_downstream_read_data_valid_sdram_s1),
      .std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register (std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register),
      .std_2s60_burst_15_downstream_requests_sdram_s1                       (std_2s60_burst_15_downstream_requests_sdram_s1),
      .std_2s60_burst_15_downstream_write                                   (std_2s60_burst_15_downstream_write),
      .std_2s60_burst_15_downstream_writedata                               (std_2s60_burst_15_downstream_writedata),
      .std_2s60_burst_16_downstream_address_to_slave                        (std_2s60_burst_16_downstream_address_to_slave),
      .std_2s60_burst_16_downstream_arbitrationshare                        (std_2s60_burst_16_downstream_arbitrationshare),
      .std_2s60_burst_16_downstream_burstcount                              (std_2s60_burst_16_downstream_burstcount),
      .std_2s60_burst_16_downstream_byteenable                              (std_2s60_burst_16_downstream_byteenable),
      .std_2s60_burst_16_downstream_granted_sdram_s1                        (std_2s60_burst_16_downstream_granted_sdram_s1),
      .std_2s60_burst_16_downstream_latency_counter                         (std_2s60_burst_16_downstream_latency_counter),
      .std_2s60_burst_16_downstream_qualified_request_sdram_s1              (std_2s60_burst_16_downstream_qualified_request_sdram_s1),
      .std_2s60_burst_16_downstream_read                                    (std_2s60_burst_16_downstream_read),
      .std_2s60_burst_16_downstream_read_data_valid_sdram_s1                (std_2s60_burst_16_downstream_read_data_valid_sdram_s1),
      .std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register (std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register),
      .std_2s60_burst_16_downstream_requests_sdram_s1                       (std_2s60_burst_16_downstream_requests_sdram_s1),
      .std_2s60_burst_16_downstream_write                                   (std_2s60_burst_16_downstream_write),
      .std_2s60_burst_16_downstream_writedata                               (std_2s60_burst_16_downstream_writedata)
    );

  sdram the_sdram
    (
      .az_addr        (sdram_s1_address),
      .az_be_n        (sdram_s1_byteenable_n),
      .az_cs          (sdram_s1_chipselect),
      .az_data        (sdram_s1_writedata),
      .az_rd_n        (sdram_s1_read_n),
      .az_wr_n        (sdram_s1_write_n),
      .clk            (clk),
      .reset_n        (sdram_s1_reset_n),
      .za_data        (sdram_s1_readdata),
      .za_valid       (sdram_s1_readdatavalid),
      .za_waitrequest (sdram_s1_waitrequest),
      .zs_addr        (zs_addr_from_the_sdram),
      .zs_ba          (zs_ba_from_the_sdram),
      .zs_cas_n       (zs_cas_n_from_the_sdram),
      .zs_cke         (zs_cke_from_the_sdram),
      .zs_cs_n        (zs_cs_n_from_the_sdram),
      .zs_dq          (zs_dq_to_and_from_the_sdram),
      .zs_dqm         (zs_dqm_from_the_sdram),
      .zs_ras_n       (zs_ras_n_from_the_sdram),
      .zs_we_n        (zs_we_n_from_the_sdram)
    );

  std_2s60_burst_0_upstream_arbitrator the_std_2s60_burst_0_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_0_upstream                         (cpu_instruction_master_granted_std_2s60_burst_0_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_0_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_0_upstream                        (cpu_instruction_master_requests_std_2s60_burst_0_upstream),
      .d1_std_2s60_burst_0_upstream_end_xfer                                            (d1_std_2s60_burst_0_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_0_upstream_address                                                (std_2s60_burst_0_upstream_address),
      .std_2s60_burst_0_upstream_byteaddress                                            (std_2s60_burst_0_upstream_byteaddress),
      .std_2s60_burst_0_upstream_byteenable                                             (std_2s60_burst_0_upstream_byteenable),
      .std_2s60_burst_0_upstream_debugaccess                                            (std_2s60_burst_0_upstream_debugaccess),
      .std_2s60_burst_0_upstream_read                                                   (std_2s60_burst_0_upstream_read),
      .std_2s60_burst_0_upstream_readdata                                               (std_2s60_burst_0_upstream_readdata),
      .std_2s60_burst_0_upstream_readdata_from_sa                                       (std_2s60_burst_0_upstream_readdata_from_sa),
      .std_2s60_burst_0_upstream_readdatavalid                                          (std_2s60_burst_0_upstream_readdatavalid),
      .std_2s60_burst_0_upstream_waitrequest                                            (std_2s60_burst_0_upstream_waitrequest),
      .std_2s60_burst_0_upstream_waitrequest_from_sa                                    (std_2s60_burst_0_upstream_waitrequest_from_sa),
      .std_2s60_burst_0_upstream_write                                                  (std_2s60_burst_0_upstream_write)
    );

  std_2s60_burst_0_downstream_arbitrator the_std_2s60_burst_0_downstream
    (
      .clk                                                                 (clk),
      .cpu_jtag_debug_module_readdata_from_sa                              (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                                   (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                             (clk_reset_n),
      .std_2s60_burst_0_downstream_address                                 (std_2s60_burst_0_downstream_address),
      .std_2s60_burst_0_downstream_address_to_slave                        (std_2s60_burst_0_downstream_address_to_slave),
      .std_2s60_burst_0_downstream_burstcount                              (std_2s60_burst_0_downstream_burstcount),
      .std_2s60_burst_0_downstream_byteenable                              (std_2s60_burst_0_downstream_byteenable),
      .std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module           (std_2s60_burst_0_downstream_granted_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_latency_counter                         (std_2s60_burst_0_downstream_latency_counter),
      .std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module (std_2s60_burst_0_downstream_qualified_request_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_read                                    (std_2s60_burst_0_downstream_read),
      .std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module   (std_2s60_burst_0_downstream_read_data_valid_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_readdata                                (std_2s60_burst_0_downstream_readdata),
      .std_2s60_burst_0_downstream_readdatavalid                           (std_2s60_burst_0_downstream_readdatavalid),
      .std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module          (std_2s60_burst_0_downstream_requests_cpu_jtag_debug_module),
      .std_2s60_burst_0_downstream_reset_n                                 (std_2s60_burst_0_downstream_reset_n),
      .std_2s60_burst_0_downstream_waitrequest                             (std_2s60_burst_0_downstream_waitrequest),
      .std_2s60_burst_0_downstream_write                                   (std_2s60_burst_0_downstream_write),
      .std_2s60_burst_0_downstream_writedata                               (std_2s60_burst_0_downstream_writedata)
    );

  std_2s60_burst_0 the_std_2s60_burst_0
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_0_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_0_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_0_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_0_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_0_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_0_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_0_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_0_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_0_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_0_downstream_read),
      .reg_downstream_write            (std_2s60_burst_0_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_0_downstream_writedata),
      .reset_n                         (std_2s60_burst_0_downstream_reset_n),
      .upstream_address                (std_2s60_burst_0_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_0_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_0_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_0_upstream_address),
      .upstream_read                   (std_2s60_burst_0_upstream_read),
      .upstream_readdata               (std_2s60_burst_0_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_0_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_0_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_0_upstream_write),
      .upstream_writedata              (std_2s60_burst_0_upstream_writedata)
    );

  std_2s60_burst_1_upstream_arbitrator the_std_2s60_burst_1_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_1_upstream                         (cpu_data_master_granted_std_2s60_burst_1_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_1_upstream               (cpu_data_master_qualified_request_std_2s60_burst_1_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_1_upstream                        (cpu_data_master_requests_std_2s60_burst_1_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_1_upstream_end_xfer                                     (d1_std_2s60_burst_1_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_1_upstream_address                                         (std_2s60_burst_1_upstream_address),
      .std_2s60_burst_1_upstream_burstcount                                      (std_2s60_burst_1_upstream_burstcount),
      .std_2s60_burst_1_upstream_byteaddress                                     (std_2s60_burst_1_upstream_byteaddress),
      .std_2s60_burst_1_upstream_byteenable                                      (std_2s60_burst_1_upstream_byteenable),
      .std_2s60_burst_1_upstream_debugaccess                                     (std_2s60_burst_1_upstream_debugaccess),
      .std_2s60_burst_1_upstream_read                                            (std_2s60_burst_1_upstream_read),
      .std_2s60_burst_1_upstream_readdata                                        (std_2s60_burst_1_upstream_readdata),
      .std_2s60_burst_1_upstream_readdata_from_sa                                (std_2s60_burst_1_upstream_readdata_from_sa),
      .std_2s60_burst_1_upstream_readdatavalid                                   (std_2s60_burst_1_upstream_readdatavalid),
      .std_2s60_burst_1_upstream_waitrequest                                     (std_2s60_burst_1_upstream_waitrequest),
      .std_2s60_burst_1_upstream_waitrequest_from_sa                             (std_2s60_burst_1_upstream_waitrequest_from_sa),
      .std_2s60_burst_1_upstream_write                                           (std_2s60_burst_1_upstream_write),
      .std_2s60_burst_1_upstream_writedata                                       (std_2s60_burst_1_upstream_writedata)
    );

  std_2s60_burst_1_downstream_arbitrator the_std_2s60_burst_1_downstream
    (
      .clk                                                                 (clk),
      .cpu_jtag_debug_module_readdata_from_sa                              (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                                   (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                             (clk_reset_n),
      .std_2s60_burst_1_downstream_address                                 (std_2s60_burst_1_downstream_address),
      .std_2s60_burst_1_downstream_address_to_slave                        (std_2s60_burst_1_downstream_address_to_slave),
      .std_2s60_burst_1_downstream_burstcount                              (std_2s60_burst_1_downstream_burstcount),
      .std_2s60_burst_1_downstream_byteenable                              (std_2s60_burst_1_downstream_byteenable),
      .std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module           (std_2s60_burst_1_downstream_granted_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_latency_counter                         (std_2s60_burst_1_downstream_latency_counter),
      .std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module (std_2s60_burst_1_downstream_qualified_request_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_read                                    (std_2s60_burst_1_downstream_read),
      .std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module   (std_2s60_burst_1_downstream_read_data_valid_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_readdata                                (std_2s60_burst_1_downstream_readdata),
      .std_2s60_burst_1_downstream_readdatavalid                           (std_2s60_burst_1_downstream_readdatavalid),
      .std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module          (std_2s60_burst_1_downstream_requests_cpu_jtag_debug_module),
      .std_2s60_burst_1_downstream_reset_n                                 (std_2s60_burst_1_downstream_reset_n),
      .std_2s60_burst_1_downstream_waitrequest                             (std_2s60_burst_1_downstream_waitrequest),
      .std_2s60_burst_1_downstream_write                                   (std_2s60_burst_1_downstream_write),
      .std_2s60_burst_1_downstream_writedata                               (std_2s60_burst_1_downstream_writedata)
    );

  std_2s60_burst_1 the_std_2s60_burst_1
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_1_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_1_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_1_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_1_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_1_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_1_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_1_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_1_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_1_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_1_downstream_read),
      .reg_downstream_write            (std_2s60_burst_1_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_1_downstream_writedata),
      .reset_n                         (std_2s60_burst_1_downstream_reset_n),
      .upstream_address                (std_2s60_burst_1_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_1_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_1_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_1_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_1_upstream_address),
      .upstream_read                   (std_2s60_burst_1_upstream_read),
      .upstream_readdata               (std_2s60_burst_1_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_1_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_1_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_1_upstream_write),
      .upstream_writedata              (std_2s60_burst_1_upstream_writedata)
    );

  std_2s60_burst_10_upstream_arbitrator the_std_2s60_burst_10_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_10_upstream                        (cpu_data_master_granted_std_2s60_burst_10_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_10_upstream              (cpu_data_master_qualified_request_std_2s60_burst_10_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_10_upstream                       (cpu_data_master_requests_std_2s60_burst_10_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_10_upstream_end_xfer                                    (d1_std_2s60_burst_10_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_10_upstream_address                                        (std_2s60_burst_10_upstream_address),
      .std_2s60_burst_10_upstream_burstcount                                     (std_2s60_burst_10_upstream_burstcount),
      .std_2s60_burst_10_upstream_byteaddress                                    (std_2s60_burst_10_upstream_byteaddress),
      .std_2s60_burst_10_upstream_byteenable                                     (std_2s60_burst_10_upstream_byteenable),
      .std_2s60_burst_10_upstream_debugaccess                                    (std_2s60_burst_10_upstream_debugaccess),
      .std_2s60_burst_10_upstream_read                                           (std_2s60_burst_10_upstream_read),
      .std_2s60_burst_10_upstream_readdata                                       (std_2s60_burst_10_upstream_readdata),
      .std_2s60_burst_10_upstream_readdata_from_sa                               (std_2s60_burst_10_upstream_readdata_from_sa),
      .std_2s60_burst_10_upstream_readdatavalid                                  (std_2s60_burst_10_upstream_readdatavalid),
      .std_2s60_burst_10_upstream_waitrequest                                    (std_2s60_burst_10_upstream_waitrequest),
      .std_2s60_burst_10_upstream_waitrequest_from_sa                            (std_2s60_burst_10_upstream_waitrequest_from_sa),
      .std_2s60_burst_10_upstream_write                                          (std_2s60_burst_10_upstream_write),
      .std_2s60_burst_10_upstream_writedata                                      (std_2s60_burst_10_upstream_writedata)
    );

  std_2s60_burst_10_downstream_arbitrator the_std_2s60_burst_10_downstream
    (
      .clk                                                             (clk),
      .d1_sys_clk_timer_s1_end_xfer                                    (d1_sys_clk_timer_s1_end_xfer),
      .reset_n                                                         (clk_reset_n),
      .std_2s60_burst_10_downstream_address                            (std_2s60_burst_10_downstream_address),
      .std_2s60_burst_10_downstream_address_to_slave                   (std_2s60_burst_10_downstream_address_to_slave),
      .std_2s60_burst_10_downstream_burstcount                         (std_2s60_burst_10_downstream_burstcount),
      .std_2s60_burst_10_downstream_byteenable                         (std_2s60_burst_10_downstream_byteenable),
      .std_2s60_burst_10_downstream_granted_sys_clk_timer_s1           (std_2s60_burst_10_downstream_granted_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_latency_counter                    (std_2s60_burst_10_downstream_latency_counter),
      .std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 (std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_read                               (std_2s60_burst_10_downstream_read),
      .std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1   (std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_readdata                           (std_2s60_burst_10_downstream_readdata),
      .std_2s60_burst_10_downstream_readdatavalid                      (std_2s60_burst_10_downstream_readdatavalid),
      .std_2s60_burst_10_downstream_requests_sys_clk_timer_s1          (std_2s60_burst_10_downstream_requests_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_reset_n                            (std_2s60_burst_10_downstream_reset_n),
      .std_2s60_burst_10_downstream_waitrequest                        (std_2s60_burst_10_downstream_waitrequest),
      .std_2s60_burst_10_downstream_write                              (std_2s60_burst_10_downstream_write),
      .std_2s60_burst_10_downstream_writedata                          (std_2s60_burst_10_downstream_writedata),
      .sys_clk_timer_s1_readdata_from_sa                               (sys_clk_timer_s1_readdata_from_sa)
    );

  std_2s60_burst_10 the_std_2s60_burst_10
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_10_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_10_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_10_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_10_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_10_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_10_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_10_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_10_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_10_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_10_downstream_read),
      .reg_downstream_write            (std_2s60_burst_10_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_10_downstream_writedata),
      .reset_n                         (std_2s60_burst_10_downstream_reset_n),
      .upstream_address                (std_2s60_burst_10_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_10_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_10_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_10_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_10_upstream_address),
      .upstream_read                   (std_2s60_burst_10_upstream_read),
      .upstream_readdata               (std_2s60_burst_10_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_10_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_10_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_10_upstream_write),
      .upstream_writedata              (std_2s60_burst_10_upstream_writedata)
    );

  std_2s60_burst_11_upstream_arbitrator the_std_2s60_burst_11_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_11_upstream                        (cpu_data_master_granted_std_2s60_burst_11_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_11_upstream              (cpu_data_master_qualified_request_std_2s60_burst_11_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_11_upstream                       (cpu_data_master_requests_std_2s60_burst_11_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_11_upstream_end_xfer                                    (d1_std_2s60_burst_11_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_11_upstream_address                                        (std_2s60_burst_11_upstream_address),
      .std_2s60_burst_11_upstream_burstcount                                     (std_2s60_burst_11_upstream_burstcount),
      .std_2s60_burst_11_upstream_byteaddress                                    (std_2s60_burst_11_upstream_byteaddress),
      .std_2s60_burst_11_upstream_byteenable                                     (std_2s60_burst_11_upstream_byteenable),
      .std_2s60_burst_11_upstream_debugaccess                                    (std_2s60_burst_11_upstream_debugaccess),
      .std_2s60_burst_11_upstream_read                                           (std_2s60_burst_11_upstream_read),
      .std_2s60_burst_11_upstream_readdata                                       (std_2s60_burst_11_upstream_readdata),
      .std_2s60_burst_11_upstream_readdata_from_sa                               (std_2s60_burst_11_upstream_readdata_from_sa),
      .std_2s60_burst_11_upstream_readdatavalid                                  (std_2s60_burst_11_upstream_readdatavalid),
      .std_2s60_burst_11_upstream_waitrequest                                    (std_2s60_burst_11_upstream_waitrequest),
      .std_2s60_burst_11_upstream_waitrequest_from_sa                            (std_2s60_burst_11_upstream_waitrequest_from_sa),
      .std_2s60_burst_11_upstream_write                                          (std_2s60_burst_11_upstream_write),
      .std_2s60_burst_11_upstream_writedata                                      (std_2s60_burst_11_upstream_writedata)
    );

  std_2s60_burst_11_downstream_arbitrator the_std_2s60_burst_11_downstream
    (
      .clk                                                                        (clk),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                    (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                               (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                            (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .reset_n                                                                    (clk_reset_n),
      .std_2s60_burst_11_downstream_address                                       (std_2s60_burst_11_downstream_address),
      .std_2s60_burst_11_downstream_address_to_slave                              (std_2s60_burst_11_downstream_address_to_slave),
      .std_2s60_burst_11_downstream_burstcount                                    (std_2s60_burst_11_downstream_burstcount),
      .std_2s60_burst_11_downstream_byteenable                                    (std_2s60_burst_11_downstream_byteenable),
      .std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave           (std_2s60_burst_11_downstream_granted_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_latency_counter                               (std_2s60_burst_11_downstream_latency_counter),
      .std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave (std_2s60_burst_11_downstream_qualified_request_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_read                                          (std_2s60_burst_11_downstream_read),
      .std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave   (std_2s60_burst_11_downstream_read_data_valid_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_readdata                                      (std_2s60_burst_11_downstream_readdata),
      .std_2s60_burst_11_downstream_readdatavalid                                 (std_2s60_burst_11_downstream_readdatavalid),
      .std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave          (std_2s60_burst_11_downstream_requests_jtag_uart_avalon_jtag_slave),
      .std_2s60_burst_11_downstream_reset_n                                       (std_2s60_burst_11_downstream_reset_n),
      .std_2s60_burst_11_downstream_waitrequest                                   (std_2s60_burst_11_downstream_waitrequest),
      .std_2s60_burst_11_downstream_write                                         (std_2s60_burst_11_downstream_write),
      .std_2s60_burst_11_downstream_writedata                                     (std_2s60_burst_11_downstream_writedata)
    );

  std_2s60_burst_11 the_std_2s60_burst_11
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_11_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_11_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_11_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_11_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_11_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_11_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_11_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_11_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_11_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_11_downstream_read),
      .reg_downstream_write            (std_2s60_burst_11_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_11_downstream_writedata),
      .reset_n                         (std_2s60_burst_11_downstream_reset_n),
      .upstream_address                (std_2s60_burst_11_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_11_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_11_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_11_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_11_upstream_address),
      .upstream_read                   (std_2s60_burst_11_upstream_read),
      .upstream_readdata               (std_2s60_burst_11_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_11_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_11_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_11_upstream_write),
      .upstream_writedata              (std_2s60_burst_11_upstream_writedata)
    );

  std_2s60_burst_12_upstream_arbitrator the_std_2s60_burst_12_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_12_upstream                        (cpu_data_master_granted_std_2s60_burst_12_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_12_upstream              (cpu_data_master_qualified_request_std_2s60_burst_12_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_12_upstream                       (cpu_data_master_requests_std_2s60_burst_12_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_12_upstream_end_xfer                                    (d1_std_2s60_burst_12_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_12_upstream_address                                        (std_2s60_burst_12_upstream_address),
      .std_2s60_burst_12_upstream_burstcount                                     (std_2s60_burst_12_upstream_burstcount),
      .std_2s60_burst_12_upstream_byteaddress                                    (std_2s60_burst_12_upstream_byteaddress),
      .std_2s60_burst_12_upstream_byteenable                                     (std_2s60_burst_12_upstream_byteenable),
      .std_2s60_burst_12_upstream_debugaccess                                    (std_2s60_burst_12_upstream_debugaccess),
      .std_2s60_burst_12_upstream_read                                           (std_2s60_burst_12_upstream_read),
      .std_2s60_burst_12_upstream_readdata                                       (std_2s60_burst_12_upstream_readdata),
      .std_2s60_burst_12_upstream_readdata_from_sa                               (std_2s60_burst_12_upstream_readdata_from_sa),
      .std_2s60_burst_12_upstream_readdatavalid                                  (std_2s60_burst_12_upstream_readdatavalid),
      .std_2s60_burst_12_upstream_waitrequest                                    (std_2s60_burst_12_upstream_waitrequest),
      .std_2s60_burst_12_upstream_waitrequest_from_sa                            (std_2s60_burst_12_upstream_waitrequest_from_sa),
      .std_2s60_burst_12_upstream_write                                          (std_2s60_burst_12_upstream_write),
      .std_2s60_burst_12_upstream_writedata                                      (std_2s60_burst_12_upstream_writedata)
    );

  std_2s60_burst_12_downstream_arbitrator the_std_2s60_burst_12_downstream
    (
      .clk                                                              (clk),
      .d1_high_res_timer_s1_end_xfer                                    (d1_high_res_timer_s1_end_xfer),
      .high_res_timer_s1_readdata_from_sa                               (high_res_timer_s1_readdata_from_sa),
      .reset_n                                                          (clk_reset_n),
      .std_2s60_burst_12_downstream_address                             (std_2s60_burst_12_downstream_address),
      .std_2s60_burst_12_downstream_address_to_slave                    (std_2s60_burst_12_downstream_address_to_slave),
      .std_2s60_burst_12_downstream_burstcount                          (std_2s60_burst_12_downstream_burstcount),
      .std_2s60_burst_12_downstream_byteenable                          (std_2s60_burst_12_downstream_byteenable),
      .std_2s60_burst_12_downstream_granted_high_res_timer_s1           (std_2s60_burst_12_downstream_granted_high_res_timer_s1),
      .std_2s60_burst_12_downstream_latency_counter                     (std_2s60_burst_12_downstream_latency_counter),
      .std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1 (std_2s60_burst_12_downstream_qualified_request_high_res_timer_s1),
      .std_2s60_burst_12_downstream_read                                (std_2s60_burst_12_downstream_read),
      .std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1   (std_2s60_burst_12_downstream_read_data_valid_high_res_timer_s1),
      .std_2s60_burst_12_downstream_readdata                            (std_2s60_burst_12_downstream_readdata),
      .std_2s60_burst_12_downstream_readdatavalid                       (std_2s60_burst_12_downstream_readdatavalid),
      .std_2s60_burst_12_downstream_requests_high_res_timer_s1          (std_2s60_burst_12_downstream_requests_high_res_timer_s1),
      .std_2s60_burst_12_downstream_reset_n                             (std_2s60_burst_12_downstream_reset_n),
      .std_2s60_burst_12_downstream_waitrequest                         (std_2s60_burst_12_downstream_waitrequest),
      .std_2s60_burst_12_downstream_write                               (std_2s60_burst_12_downstream_write),
      .std_2s60_burst_12_downstream_writedata                           (std_2s60_burst_12_downstream_writedata)
    );

  std_2s60_burst_12 the_std_2s60_burst_12
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_12_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_12_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_12_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_12_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_12_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_12_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_12_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_12_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_12_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_12_downstream_read),
      .reg_downstream_write            (std_2s60_burst_12_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_12_downstream_writedata),
      .reset_n                         (std_2s60_burst_12_downstream_reset_n),
      .upstream_address                (std_2s60_burst_12_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_12_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_12_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_12_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_12_upstream_address),
      .upstream_read                   (std_2s60_burst_12_upstream_read),
      .upstream_readdata               (std_2s60_burst_12_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_12_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_12_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_12_upstream_write),
      .upstream_writedata              (std_2s60_burst_12_upstream_writedata)
    );

  std_2s60_burst_13_upstream_arbitrator the_std_2s60_burst_13_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_13_upstream                        (cpu_data_master_granted_std_2s60_burst_13_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_13_upstream              (cpu_data_master_qualified_request_std_2s60_burst_13_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_13_upstream                       (cpu_data_master_requests_std_2s60_burst_13_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_13_upstream_end_xfer                                    (d1_std_2s60_burst_13_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_13_upstream_address                                        (std_2s60_burst_13_upstream_address),
      .std_2s60_burst_13_upstream_burstcount                                     (std_2s60_burst_13_upstream_burstcount),
      .std_2s60_burst_13_upstream_byteaddress                                    (std_2s60_burst_13_upstream_byteaddress),
      .std_2s60_burst_13_upstream_byteenable                                     (std_2s60_burst_13_upstream_byteenable),
      .std_2s60_burst_13_upstream_debugaccess                                    (std_2s60_burst_13_upstream_debugaccess),
      .std_2s60_burst_13_upstream_read                                           (std_2s60_burst_13_upstream_read),
      .std_2s60_burst_13_upstream_readdata                                       (std_2s60_burst_13_upstream_readdata),
      .std_2s60_burst_13_upstream_readdata_from_sa                               (std_2s60_burst_13_upstream_readdata_from_sa),
      .std_2s60_burst_13_upstream_readdatavalid                                  (std_2s60_burst_13_upstream_readdatavalid),
      .std_2s60_burst_13_upstream_waitrequest                                    (std_2s60_burst_13_upstream_waitrequest),
      .std_2s60_burst_13_upstream_waitrequest_from_sa                            (std_2s60_burst_13_upstream_waitrequest_from_sa),
      .std_2s60_burst_13_upstream_write                                          (std_2s60_burst_13_upstream_write),
      .std_2s60_burst_13_upstream_writedata                                      (std_2s60_burst_13_upstream_writedata)
    );

  std_2s60_burst_13_downstream_arbitrator the_std_2s60_burst_13_downstream
    (
      .clk                                                                    (clk),
      .d1_reconfig_request_pio_s1_end_xfer                                    (d1_reconfig_request_pio_s1_end_xfer),
      .reconfig_request_pio_s1_readdata_from_sa                               (reconfig_request_pio_s1_readdata_from_sa),
      .reset_n                                                                (clk_reset_n),
      .std_2s60_burst_13_downstream_address                                   (std_2s60_burst_13_downstream_address),
      .std_2s60_burst_13_downstream_address_to_slave                          (std_2s60_burst_13_downstream_address_to_slave),
      .std_2s60_burst_13_downstream_burstcount                                (std_2s60_burst_13_downstream_burstcount),
      .std_2s60_burst_13_downstream_byteenable                                (std_2s60_burst_13_downstream_byteenable),
      .std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1           (std_2s60_burst_13_downstream_granted_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_latency_counter                           (std_2s60_burst_13_downstream_latency_counter),
      .std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1 (std_2s60_burst_13_downstream_qualified_request_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_read                                      (std_2s60_burst_13_downstream_read),
      .std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1   (std_2s60_burst_13_downstream_read_data_valid_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_readdata                                  (std_2s60_burst_13_downstream_readdata),
      .std_2s60_burst_13_downstream_readdatavalid                             (std_2s60_burst_13_downstream_readdatavalid),
      .std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1          (std_2s60_burst_13_downstream_requests_reconfig_request_pio_s1),
      .std_2s60_burst_13_downstream_reset_n                                   (std_2s60_burst_13_downstream_reset_n),
      .std_2s60_burst_13_downstream_waitrequest                               (std_2s60_burst_13_downstream_waitrequest),
      .std_2s60_burst_13_downstream_write                                     (std_2s60_burst_13_downstream_write),
      .std_2s60_burst_13_downstream_writedata                                 (std_2s60_burst_13_downstream_writedata)
    );

  std_2s60_burst_13 the_std_2s60_burst_13
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_13_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_13_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_13_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_13_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_13_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_13_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_13_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_13_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_13_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_13_downstream_read),
      .reg_downstream_write            (std_2s60_burst_13_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_13_downstream_writedata),
      .reset_n                         (std_2s60_burst_13_downstream_reset_n),
      .upstream_address                (std_2s60_burst_13_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_13_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_13_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_13_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_13_upstream_address),
      .upstream_read                   (std_2s60_burst_13_upstream_read),
      .upstream_readdata               (std_2s60_burst_13_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_13_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_13_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_13_upstream_write),
      .upstream_writedata              (std_2s60_burst_13_upstream_writedata)
    );

  std_2s60_burst_14_upstream_arbitrator the_std_2s60_burst_14_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_14_upstream                        (cpu_data_master_granted_std_2s60_burst_14_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_14_upstream              (cpu_data_master_qualified_request_std_2s60_burst_14_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_14_upstream                       (cpu_data_master_requests_std_2s60_burst_14_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_14_upstream_end_xfer                                    (d1_std_2s60_burst_14_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_14_upstream_address                                        (std_2s60_burst_14_upstream_address),
      .std_2s60_burst_14_upstream_burstcount                                     (std_2s60_burst_14_upstream_burstcount),
      .std_2s60_burst_14_upstream_byteaddress                                    (std_2s60_burst_14_upstream_byteaddress),
      .std_2s60_burst_14_upstream_byteenable                                     (std_2s60_burst_14_upstream_byteenable),
      .std_2s60_burst_14_upstream_debugaccess                                    (std_2s60_burst_14_upstream_debugaccess),
      .std_2s60_burst_14_upstream_read                                           (std_2s60_burst_14_upstream_read),
      .std_2s60_burst_14_upstream_readdata                                       (std_2s60_burst_14_upstream_readdata),
      .std_2s60_burst_14_upstream_readdata_from_sa                               (std_2s60_burst_14_upstream_readdata_from_sa),
      .std_2s60_burst_14_upstream_readdatavalid                                  (std_2s60_burst_14_upstream_readdatavalid),
      .std_2s60_burst_14_upstream_waitrequest                                    (std_2s60_burst_14_upstream_waitrequest),
      .std_2s60_burst_14_upstream_waitrequest_from_sa                            (std_2s60_burst_14_upstream_waitrequest_from_sa),
      .std_2s60_burst_14_upstream_write                                          (std_2s60_burst_14_upstream_write),
      .std_2s60_burst_14_upstream_writedata                                      (std_2s60_burst_14_upstream_writedata)
    );

  std_2s60_burst_14_downstream_arbitrator the_std_2s60_burst_14_downstream
    (
      .clk                                                                (clk),
      .d1_sysid_control_slave_end_xfer                                    (d1_sysid_control_slave_end_xfer),
      .reset_n                                                            (clk_reset_n),
      .std_2s60_burst_14_downstream_address                               (std_2s60_burst_14_downstream_address),
      .std_2s60_burst_14_downstream_address_to_slave                      (std_2s60_burst_14_downstream_address_to_slave),
      .std_2s60_burst_14_downstream_burstcount                            (std_2s60_burst_14_downstream_burstcount),
      .std_2s60_burst_14_downstream_byteenable                            (std_2s60_burst_14_downstream_byteenable),
      .std_2s60_burst_14_downstream_granted_sysid_control_slave           (std_2s60_burst_14_downstream_granted_sysid_control_slave),
      .std_2s60_burst_14_downstream_latency_counter                       (std_2s60_burst_14_downstream_latency_counter),
      .std_2s60_burst_14_downstream_qualified_request_sysid_control_slave (std_2s60_burst_14_downstream_qualified_request_sysid_control_slave),
      .std_2s60_burst_14_downstream_read                                  (std_2s60_burst_14_downstream_read),
      .std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave   (std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave),
      .std_2s60_burst_14_downstream_readdata                              (std_2s60_burst_14_downstream_readdata),
      .std_2s60_burst_14_downstream_readdatavalid                         (std_2s60_burst_14_downstream_readdatavalid),
      .std_2s60_burst_14_downstream_requests_sysid_control_slave          (std_2s60_burst_14_downstream_requests_sysid_control_slave),
      .std_2s60_burst_14_downstream_reset_n                               (std_2s60_burst_14_downstream_reset_n),
      .std_2s60_burst_14_downstream_waitrequest                           (std_2s60_burst_14_downstream_waitrequest),
      .std_2s60_burst_14_downstream_write                                 (std_2s60_burst_14_downstream_write),
      .std_2s60_burst_14_downstream_writedata                             (std_2s60_burst_14_downstream_writedata),
      .sysid_control_slave_readdata_from_sa                               (sysid_control_slave_readdata_from_sa)
    );

  std_2s60_burst_14 the_std_2s60_burst_14
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_14_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_14_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_14_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_14_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_14_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_14_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_14_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_14_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_14_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_14_downstream_read),
      .reg_downstream_write            (std_2s60_burst_14_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_14_downstream_writedata),
      .reset_n                         (std_2s60_burst_14_downstream_reset_n),
      .upstream_address                (std_2s60_burst_14_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_14_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_14_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_14_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_14_upstream_address),
      .upstream_read                   (std_2s60_burst_14_upstream_read),
      .upstream_readdata               (std_2s60_burst_14_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_14_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_14_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_14_upstream_write),
      .upstream_writedata              (std_2s60_burst_14_upstream_writedata)
    );

  std_2s60_burst_15_upstream_arbitrator the_std_2s60_burst_15_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_15_upstream                        (cpu_instruction_master_granted_std_2s60_burst_15_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream              (cpu_instruction_master_qualified_request_std_2s60_burst_15_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream                (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_15_upstream                       (cpu_instruction_master_requests_std_2s60_burst_15_upstream),
      .d1_std_2s60_burst_15_upstream_end_xfer                                           (d1_std_2s60_burst_15_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_15_upstream_address                                               (std_2s60_burst_15_upstream_address),
      .std_2s60_burst_15_upstream_byteaddress                                           (std_2s60_burst_15_upstream_byteaddress),
      .std_2s60_burst_15_upstream_byteenable                                            (std_2s60_burst_15_upstream_byteenable),
      .std_2s60_burst_15_upstream_debugaccess                                           (std_2s60_burst_15_upstream_debugaccess),
      .std_2s60_burst_15_upstream_read                                                  (std_2s60_burst_15_upstream_read),
      .std_2s60_burst_15_upstream_readdata                                              (std_2s60_burst_15_upstream_readdata),
      .std_2s60_burst_15_upstream_readdata_from_sa                                      (std_2s60_burst_15_upstream_readdata_from_sa),
      .std_2s60_burst_15_upstream_readdatavalid                                         (std_2s60_burst_15_upstream_readdatavalid),
      .std_2s60_burst_15_upstream_waitrequest                                           (std_2s60_burst_15_upstream_waitrequest),
      .std_2s60_burst_15_upstream_waitrequest_from_sa                                   (std_2s60_burst_15_upstream_waitrequest_from_sa),
      .std_2s60_burst_15_upstream_write                                                 (std_2s60_burst_15_upstream_write)
    );

  std_2s60_burst_15_downstream_arbitrator the_std_2s60_burst_15_downstream
    (
      .clk                                                                  (clk),
      .d1_sdram_s1_end_xfer                                                 (d1_sdram_s1_end_xfer),
      .reset_n                                                              (clk_reset_n),
      .sdram_s1_readdata_from_sa                                            (sdram_s1_readdata_from_sa),
      .sdram_s1_waitrequest_from_sa                                         (sdram_s1_waitrequest_from_sa),
      .std_2s60_burst_15_downstream_address                                 (std_2s60_burst_15_downstream_address),
      .std_2s60_burst_15_downstream_address_to_slave                        (std_2s60_burst_15_downstream_address_to_slave),
      .std_2s60_burst_15_downstream_burstcount                              (std_2s60_burst_15_downstream_burstcount),
      .std_2s60_burst_15_downstream_byteenable                              (std_2s60_burst_15_downstream_byteenable),
      .std_2s60_burst_15_downstream_granted_sdram_s1                        (std_2s60_burst_15_downstream_granted_sdram_s1),
      .std_2s60_burst_15_downstream_latency_counter                         (std_2s60_burst_15_downstream_latency_counter),
      .std_2s60_burst_15_downstream_qualified_request_sdram_s1              (std_2s60_burst_15_downstream_qualified_request_sdram_s1),
      .std_2s60_burst_15_downstream_read                                    (std_2s60_burst_15_downstream_read),
      .std_2s60_burst_15_downstream_read_data_valid_sdram_s1                (std_2s60_burst_15_downstream_read_data_valid_sdram_s1),
      .std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register (std_2s60_burst_15_downstream_read_data_valid_sdram_s1_shift_register),
      .std_2s60_burst_15_downstream_readdata                                (std_2s60_burst_15_downstream_readdata),
      .std_2s60_burst_15_downstream_readdatavalid                           (std_2s60_burst_15_downstream_readdatavalid),
      .std_2s60_burst_15_downstream_requests_sdram_s1                       (std_2s60_burst_15_downstream_requests_sdram_s1),
      .std_2s60_burst_15_downstream_reset_n                                 (std_2s60_burst_15_downstream_reset_n),
      .std_2s60_burst_15_downstream_waitrequest                             (std_2s60_burst_15_downstream_waitrequest),
      .std_2s60_burst_15_downstream_write                                   (std_2s60_burst_15_downstream_write),
      .std_2s60_burst_15_downstream_writedata                               (std_2s60_burst_15_downstream_writedata)
    );

  std_2s60_burst_15 the_std_2s60_burst_15
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_15_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_15_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_15_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_15_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_15_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_15_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_15_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_15_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_15_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_15_downstream_read),
      .reg_downstream_write            (std_2s60_burst_15_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_15_downstream_writedata),
      .reset_n                         (std_2s60_burst_15_downstream_reset_n),
      .upstream_address                (std_2s60_burst_15_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_15_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_15_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_15_upstream_address),
      .upstream_read                   (std_2s60_burst_15_upstream_read),
      .upstream_readdata               (std_2s60_burst_15_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_15_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_15_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_15_upstream_write),
      .upstream_writedata              (std_2s60_burst_15_upstream_writedata)
    );

  std_2s60_burst_16_upstream_arbitrator the_std_2s60_burst_16_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_16_upstream                        (cpu_data_master_granted_std_2s60_burst_16_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_16_upstream              (cpu_data_master_qualified_request_std_2s60_burst_16_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_16_upstream                       (cpu_data_master_requests_std_2s60_burst_16_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_16_upstream_end_xfer                                    (d1_std_2s60_burst_16_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_16_upstream_address                                        (std_2s60_burst_16_upstream_address),
      .std_2s60_burst_16_upstream_burstcount                                     (std_2s60_burst_16_upstream_burstcount),
      .std_2s60_burst_16_upstream_byteaddress                                    (std_2s60_burst_16_upstream_byteaddress),
      .std_2s60_burst_16_upstream_byteenable                                     (std_2s60_burst_16_upstream_byteenable),
      .std_2s60_burst_16_upstream_debugaccess                                    (std_2s60_burst_16_upstream_debugaccess),
      .std_2s60_burst_16_upstream_read                                           (std_2s60_burst_16_upstream_read),
      .std_2s60_burst_16_upstream_readdata                                       (std_2s60_burst_16_upstream_readdata),
      .std_2s60_burst_16_upstream_readdata_from_sa                               (std_2s60_burst_16_upstream_readdata_from_sa),
      .std_2s60_burst_16_upstream_readdatavalid                                  (std_2s60_burst_16_upstream_readdatavalid),
      .std_2s60_burst_16_upstream_waitrequest                                    (std_2s60_burst_16_upstream_waitrequest),
      .std_2s60_burst_16_upstream_waitrequest_from_sa                            (std_2s60_burst_16_upstream_waitrequest_from_sa),
      .std_2s60_burst_16_upstream_write                                          (std_2s60_burst_16_upstream_write),
      .std_2s60_burst_16_upstream_writedata                                      (std_2s60_burst_16_upstream_writedata)
    );

  std_2s60_burst_16_downstream_arbitrator the_std_2s60_burst_16_downstream
    (
      .clk                                                                  (clk),
      .d1_sdram_s1_end_xfer                                                 (d1_sdram_s1_end_xfer),
      .reset_n                                                              (clk_reset_n),
      .sdram_s1_readdata_from_sa                                            (sdram_s1_readdata_from_sa),
      .sdram_s1_waitrequest_from_sa                                         (sdram_s1_waitrequest_from_sa),
      .std_2s60_burst_16_downstream_address                                 (std_2s60_burst_16_downstream_address),
      .std_2s60_burst_16_downstream_address_to_slave                        (std_2s60_burst_16_downstream_address_to_slave),
      .std_2s60_burst_16_downstream_burstcount                              (std_2s60_burst_16_downstream_burstcount),
      .std_2s60_burst_16_downstream_byteenable                              (std_2s60_burst_16_downstream_byteenable),
      .std_2s60_burst_16_downstream_granted_sdram_s1                        (std_2s60_burst_16_downstream_granted_sdram_s1),
      .std_2s60_burst_16_downstream_latency_counter                         (std_2s60_burst_16_downstream_latency_counter),
      .std_2s60_burst_16_downstream_qualified_request_sdram_s1              (std_2s60_burst_16_downstream_qualified_request_sdram_s1),
      .std_2s60_burst_16_downstream_read                                    (std_2s60_burst_16_downstream_read),
      .std_2s60_burst_16_downstream_read_data_valid_sdram_s1                (std_2s60_burst_16_downstream_read_data_valid_sdram_s1),
      .std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register (std_2s60_burst_16_downstream_read_data_valid_sdram_s1_shift_register),
      .std_2s60_burst_16_downstream_readdata                                (std_2s60_burst_16_downstream_readdata),
      .std_2s60_burst_16_downstream_readdatavalid                           (std_2s60_burst_16_downstream_readdatavalid),
      .std_2s60_burst_16_downstream_requests_sdram_s1                       (std_2s60_burst_16_downstream_requests_sdram_s1),
      .std_2s60_burst_16_downstream_reset_n                                 (std_2s60_burst_16_downstream_reset_n),
      .std_2s60_burst_16_downstream_waitrequest                             (std_2s60_burst_16_downstream_waitrequest),
      .std_2s60_burst_16_downstream_write                                   (std_2s60_burst_16_downstream_write),
      .std_2s60_burst_16_downstream_writedata                               (std_2s60_burst_16_downstream_writedata)
    );

  std_2s60_burst_16 the_std_2s60_burst_16
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_16_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_16_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_16_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_16_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_16_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_16_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_16_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_16_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_16_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_16_downstream_read),
      .reg_downstream_write            (std_2s60_burst_16_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_16_downstream_writedata),
      .reset_n                         (std_2s60_burst_16_downstream_reset_n),
      .upstream_address                (std_2s60_burst_16_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_16_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_16_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_16_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_16_upstream_address),
      .upstream_read                   (std_2s60_burst_16_upstream_read),
      .upstream_readdata               (std_2s60_burst_16_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_16_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_16_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_16_upstream_write),
      .upstream_writedata              (std_2s60_burst_16_upstream_writedata)
    );

  std_2s60_burst_17_upstream_arbitrator the_std_2s60_burst_17_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_17_upstream                        (cpu_data_master_granted_std_2s60_burst_17_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_17_upstream              (cpu_data_master_qualified_request_std_2s60_burst_17_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream                (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_17_upstream                       (cpu_data_master_requests_std_2s60_burst_17_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_17_upstream_end_xfer                                    (d1_std_2s60_burst_17_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_17_upstream_address                                        (std_2s60_burst_17_upstream_address),
      .std_2s60_burst_17_upstream_burstcount                                     (std_2s60_burst_17_upstream_burstcount),
      .std_2s60_burst_17_upstream_byteaddress                                    (std_2s60_burst_17_upstream_byteaddress),
      .std_2s60_burst_17_upstream_byteenable                                     (std_2s60_burst_17_upstream_byteenable),
      .std_2s60_burst_17_upstream_debugaccess                                    (std_2s60_burst_17_upstream_debugaccess),
      .std_2s60_burst_17_upstream_read                                           (std_2s60_burst_17_upstream_read),
      .std_2s60_burst_17_upstream_readdata                                       (std_2s60_burst_17_upstream_readdata),
      .std_2s60_burst_17_upstream_readdata_from_sa                               (std_2s60_burst_17_upstream_readdata_from_sa),
      .std_2s60_burst_17_upstream_readdatavalid                                  (std_2s60_burst_17_upstream_readdatavalid),
      .std_2s60_burst_17_upstream_waitrequest                                    (std_2s60_burst_17_upstream_waitrequest),
      .std_2s60_burst_17_upstream_waitrequest_from_sa                            (std_2s60_burst_17_upstream_waitrequest_from_sa),
      .std_2s60_burst_17_upstream_write                                          (std_2s60_burst_17_upstream_write),
      .std_2s60_burst_17_upstream_writedata                                      (std_2s60_burst_17_upstream_writedata)
    );

  std_2s60_burst_17_downstream_arbitrator the_std_2s60_burst_17_downstream
    (
      .ad_buf_s1_readdata_from_sa                               (ad_buf_s1_readdata_from_sa),
      .ad_buf_s1_waitrequest_from_sa                            (ad_buf_s1_waitrequest_from_sa),
      .clk                                                      (clk),
      .d1_ad_buf_s1_end_xfer                                    (d1_ad_buf_s1_end_xfer),
      .reset_n                                                  (clk_reset_n),
      .std_2s60_burst_17_downstream_address                     (std_2s60_burst_17_downstream_address),
      .std_2s60_burst_17_downstream_address_to_slave            (std_2s60_burst_17_downstream_address_to_slave),
      .std_2s60_burst_17_downstream_burstcount                  (std_2s60_burst_17_downstream_burstcount),
      .std_2s60_burst_17_downstream_byteenable                  (std_2s60_burst_17_downstream_byteenable),
      .std_2s60_burst_17_downstream_granted_ad_buf_s1           (std_2s60_burst_17_downstream_granted_ad_buf_s1),
      .std_2s60_burst_17_downstream_latency_counter             (std_2s60_burst_17_downstream_latency_counter),
      .std_2s60_burst_17_downstream_qualified_request_ad_buf_s1 (std_2s60_burst_17_downstream_qualified_request_ad_buf_s1),
      .std_2s60_burst_17_downstream_read                        (std_2s60_burst_17_downstream_read),
      .std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1   (std_2s60_burst_17_downstream_read_data_valid_ad_buf_s1),
      .std_2s60_burst_17_downstream_readdata                    (std_2s60_burst_17_downstream_readdata),
      .std_2s60_burst_17_downstream_readdatavalid               (std_2s60_burst_17_downstream_readdatavalid),
      .std_2s60_burst_17_downstream_requests_ad_buf_s1          (std_2s60_burst_17_downstream_requests_ad_buf_s1),
      .std_2s60_burst_17_downstream_reset_n                     (std_2s60_burst_17_downstream_reset_n),
      .std_2s60_burst_17_downstream_waitrequest                 (std_2s60_burst_17_downstream_waitrequest),
      .std_2s60_burst_17_downstream_write                       (std_2s60_burst_17_downstream_write),
      .std_2s60_burst_17_downstream_writedata                   (std_2s60_burst_17_downstream_writedata)
    );

  std_2s60_burst_17 the_std_2s60_burst_17
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_17_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_17_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_17_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_17_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_17_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_17_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_17_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_17_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_17_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_17_downstream_read),
      .reg_downstream_write            (std_2s60_burst_17_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_17_downstream_writedata),
      .reset_n                         (std_2s60_burst_17_downstream_reset_n),
      .upstream_address                (std_2s60_burst_17_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_17_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_17_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_17_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_17_upstream_address),
      .upstream_read                   (std_2s60_burst_17_upstream_read),
      .upstream_readdata               (std_2s60_burst_17_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_17_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_17_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_17_upstream_write),
      .upstream_writedata              (std_2s60_burst_17_upstream_writedata)
    );

  std_2s60_burst_18_upstream_arbitrator the_std_2s60_burst_18_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_18_upstream                        (cpu_instruction_master_granted_std_2s60_burst_18_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream              (cpu_instruction_master_qualified_request_std_2s60_burst_18_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream                (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_18_upstream                       (cpu_instruction_master_requests_std_2s60_burst_18_upstream),
      .d1_std_2s60_burst_18_upstream_end_xfer                                           (d1_std_2s60_burst_18_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_18_upstream_address                                               (std_2s60_burst_18_upstream_address),
      .std_2s60_burst_18_upstream_byteaddress                                           (std_2s60_burst_18_upstream_byteaddress),
      .std_2s60_burst_18_upstream_byteenable                                            (std_2s60_burst_18_upstream_byteenable),
      .std_2s60_burst_18_upstream_debugaccess                                           (std_2s60_burst_18_upstream_debugaccess),
      .std_2s60_burst_18_upstream_read                                                  (std_2s60_burst_18_upstream_read),
      .std_2s60_burst_18_upstream_readdata                                              (std_2s60_burst_18_upstream_readdata),
      .std_2s60_burst_18_upstream_readdata_from_sa                                      (std_2s60_burst_18_upstream_readdata_from_sa),
      .std_2s60_burst_18_upstream_readdatavalid                                         (std_2s60_burst_18_upstream_readdatavalid),
      .std_2s60_burst_18_upstream_waitrequest                                           (std_2s60_burst_18_upstream_waitrequest),
      .std_2s60_burst_18_upstream_waitrequest_from_sa                                   (std_2s60_burst_18_upstream_waitrequest_from_sa),
      .std_2s60_burst_18_upstream_write                                                 (std_2s60_burst_18_upstream_write)
    );

  std_2s60_burst_18_downstream_arbitrator the_std_2s60_burst_18_downstream
    (
      .ad_buf_s1_readdata_from_sa                               (ad_buf_s1_readdata_from_sa),
      .ad_buf_s1_waitrequest_from_sa                            (ad_buf_s1_waitrequest_from_sa),
      .clk                                                      (clk),
      .d1_ad_buf_s1_end_xfer                                    (d1_ad_buf_s1_end_xfer),
      .reset_n                                                  (clk_reset_n),
      .std_2s60_burst_18_downstream_address                     (std_2s60_burst_18_downstream_address),
      .std_2s60_burst_18_downstream_address_to_slave            (std_2s60_burst_18_downstream_address_to_slave),
      .std_2s60_burst_18_downstream_burstcount                  (std_2s60_burst_18_downstream_burstcount),
      .std_2s60_burst_18_downstream_byteenable                  (std_2s60_burst_18_downstream_byteenable),
      .std_2s60_burst_18_downstream_granted_ad_buf_s1           (std_2s60_burst_18_downstream_granted_ad_buf_s1),
      .std_2s60_burst_18_downstream_latency_counter             (std_2s60_burst_18_downstream_latency_counter),
      .std_2s60_burst_18_downstream_qualified_request_ad_buf_s1 (std_2s60_burst_18_downstream_qualified_request_ad_buf_s1),
      .std_2s60_burst_18_downstream_read                        (std_2s60_burst_18_downstream_read),
      .std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1   (std_2s60_burst_18_downstream_read_data_valid_ad_buf_s1),
      .std_2s60_burst_18_downstream_readdata                    (std_2s60_burst_18_downstream_readdata),
      .std_2s60_burst_18_downstream_readdatavalid               (std_2s60_burst_18_downstream_readdatavalid),
      .std_2s60_burst_18_downstream_requests_ad_buf_s1          (std_2s60_burst_18_downstream_requests_ad_buf_s1),
      .std_2s60_burst_18_downstream_reset_n                     (std_2s60_burst_18_downstream_reset_n),
      .std_2s60_burst_18_downstream_waitrequest                 (std_2s60_burst_18_downstream_waitrequest),
      .std_2s60_burst_18_downstream_write                       (std_2s60_burst_18_downstream_write),
      .std_2s60_burst_18_downstream_writedata                   (std_2s60_burst_18_downstream_writedata)
    );

  std_2s60_burst_18 the_std_2s60_burst_18
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_18_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_18_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_18_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_18_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_18_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_18_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_18_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_18_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_18_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_18_downstream_read),
      .reg_downstream_write            (std_2s60_burst_18_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_18_downstream_writedata),
      .reset_n                         (std_2s60_burst_18_downstream_reset_n),
      .upstream_address                (std_2s60_burst_18_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_18_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_18_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_18_upstream_address),
      .upstream_read                   (std_2s60_burst_18_upstream_read),
      .upstream_readdata               (std_2s60_burst_18_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_18_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_18_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_18_upstream_write),
      .upstream_writedata              (std_2s60_burst_18_upstream_writedata)
    );

  std_2s60_burst_2_upstream_arbitrator the_std_2s60_burst_2_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_dbs_address                                               (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_std_2s60_burst_2_upstream                         (cpu_instruction_master_granted_std_2s60_burst_2_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_2_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_2_upstream                        (cpu_instruction_master_requests_std_2s60_burst_2_upstream),
      .d1_std_2s60_burst_2_upstream_end_xfer                                            (d1_std_2s60_burst_2_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_2_upstream_address                                                (std_2s60_burst_2_upstream_address),
      .std_2s60_burst_2_upstream_byteaddress                                            (std_2s60_burst_2_upstream_byteaddress),
      .std_2s60_burst_2_upstream_byteenable                                             (std_2s60_burst_2_upstream_byteenable),
      .std_2s60_burst_2_upstream_debugaccess                                            (std_2s60_burst_2_upstream_debugaccess),
      .std_2s60_burst_2_upstream_read                                                   (std_2s60_burst_2_upstream_read),
      .std_2s60_burst_2_upstream_readdata                                               (std_2s60_burst_2_upstream_readdata),
      .std_2s60_burst_2_upstream_readdata_from_sa                                       (std_2s60_burst_2_upstream_readdata_from_sa),
      .std_2s60_burst_2_upstream_readdatavalid                                          (std_2s60_burst_2_upstream_readdatavalid),
      .std_2s60_burst_2_upstream_waitrequest                                            (std_2s60_burst_2_upstream_waitrequest),
      .std_2s60_burst_2_upstream_waitrequest_from_sa                                    (std_2s60_burst_2_upstream_waitrequest_from_sa),
      .std_2s60_burst_2_upstream_write                                                  (std_2s60_burst_2_upstream_write)
    );

  std_2s60_burst_2_downstream_arbitrator the_std_2s60_burst_2_downstream
    (
      .clk                                                        (clk),
      .d1_ext_flash_bus_avalon_slave_end_xfer                     (d1_ext_flash_bus_avalon_slave_end_xfer),
      .ext_flash_s1_wait_counter_eq_0                             (ext_flash_s1_wait_counter_eq_0),
      .incoming_ext_flash_bus_data_with_Xs_converted_to_0         (incoming_ext_flash_bus_data_with_Xs_converted_to_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_2_downstream_address                        (std_2s60_burst_2_downstream_address),
      .std_2s60_burst_2_downstream_address_to_slave               (std_2s60_burst_2_downstream_address_to_slave),
      .std_2s60_burst_2_downstream_burstcount                     (std_2s60_burst_2_downstream_burstcount),
      .std_2s60_burst_2_downstream_byteenable                     (std_2s60_burst_2_downstream_byteenable),
      .std_2s60_burst_2_downstream_granted_ext_flash_s1           (std_2s60_burst_2_downstream_granted_ext_flash_s1),
      .std_2s60_burst_2_downstream_latency_counter                (std_2s60_burst_2_downstream_latency_counter),
      .std_2s60_burst_2_downstream_qualified_request_ext_flash_s1 (std_2s60_burst_2_downstream_qualified_request_ext_flash_s1),
      .std_2s60_burst_2_downstream_read                           (std_2s60_burst_2_downstream_read),
      .std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1   (std_2s60_burst_2_downstream_read_data_valid_ext_flash_s1),
      .std_2s60_burst_2_downstream_readdata                       (std_2s60_burst_2_downstream_readdata),
      .std_2s60_burst_2_downstream_readdatavalid                  (std_2s60_burst_2_downstream_readdatavalid),
      .std_2s60_burst_2_downstream_requests_ext_flash_s1          (std_2s60_burst_2_downstream_requests_ext_flash_s1),
      .std_2s60_burst_2_downstream_reset_n                        (std_2s60_burst_2_downstream_reset_n),
      .std_2s60_burst_2_downstream_waitrequest                    (std_2s60_burst_2_downstream_waitrequest),
      .std_2s60_burst_2_downstream_write                          (std_2s60_burst_2_downstream_write),
      .std_2s60_burst_2_downstream_writedata                      (std_2s60_burst_2_downstream_writedata)
    );

  std_2s60_burst_2 the_std_2s60_burst_2
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_2_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_2_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_2_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_2_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_2_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_2_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_2_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_2_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_2_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_2_downstream_read),
      .reg_downstream_write            (std_2s60_burst_2_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_2_downstream_writedata),
      .reset_n                         (std_2s60_burst_2_downstream_reset_n),
      .upstream_address                (std_2s60_burst_2_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_2_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_2_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_2_upstream_address),
      .upstream_read                   (std_2s60_burst_2_upstream_read),
      .upstream_readdata               (std_2s60_burst_2_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_2_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_2_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_2_upstream_write),
      .upstream_writedata              (std_2s60_burst_2_upstream_writedata)
    );

  std_2s60_burst_3_upstream_arbitrator the_std_2s60_burst_3_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_byteenable_std_2s60_burst_3_upstream                      (cpu_data_master_byteenable_std_2s60_burst_3_upstream),
      .cpu_data_master_dbs_address                                               (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_8                                               (cpu_data_master_dbs_write_8),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_3_upstream                         (cpu_data_master_granted_std_2s60_burst_3_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_3_upstream               (cpu_data_master_qualified_request_std_2s60_burst_3_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_3_upstream                        (cpu_data_master_requests_std_2s60_burst_3_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .d1_std_2s60_burst_3_upstream_end_xfer                                     (d1_std_2s60_burst_3_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_3_upstream_address                                         (std_2s60_burst_3_upstream_address),
      .std_2s60_burst_3_upstream_burstcount                                      (std_2s60_burst_3_upstream_burstcount),
      .std_2s60_burst_3_upstream_byteaddress                                     (std_2s60_burst_3_upstream_byteaddress),
      .std_2s60_burst_3_upstream_byteenable                                      (std_2s60_burst_3_upstream_byteenable),
      .std_2s60_burst_3_upstream_debugaccess                                     (std_2s60_burst_3_upstream_debugaccess),
      .std_2s60_burst_3_upstream_read                                            (std_2s60_burst_3_upstream_read),
      .std_2s60_burst_3_upstream_readdata                                        (std_2s60_burst_3_upstream_readdata),
      .std_2s60_burst_3_upstream_readdata_from_sa                                (std_2s60_burst_3_upstream_readdata_from_sa),
      .std_2s60_burst_3_upstream_readdatavalid                                   (std_2s60_burst_3_upstream_readdatavalid),
      .std_2s60_burst_3_upstream_waitrequest                                     (std_2s60_burst_3_upstream_waitrequest),
      .std_2s60_burst_3_upstream_waitrequest_from_sa                             (std_2s60_burst_3_upstream_waitrequest_from_sa),
      .std_2s60_burst_3_upstream_write                                           (std_2s60_burst_3_upstream_write),
      .std_2s60_burst_3_upstream_writedata                                       (std_2s60_burst_3_upstream_writedata)
    );

  std_2s60_burst_3_downstream_arbitrator the_std_2s60_burst_3_downstream
    (
      .clk                                                        (clk),
      .d1_ext_flash_bus_avalon_slave_end_xfer                     (d1_ext_flash_bus_avalon_slave_end_xfer),
      .ext_flash_s1_wait_counter_eq_0                             (ext_flash_s1_wait_counter_eq_0),
      .incoming_ext_flash_bus_data_with_Xs_converted_to_0         (incoming_ext_flash_bus_data_with_Xs_converted_to_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_3_downstream_address                        (std_2s60_burst_3_downstream_address),
      .std_2s60_burst_3_downstream_address_to_slave               (std_2s60_burst_3_downstream_address_to_slave),
      .std_2s60_burst_3_downstream_burstcount                     (std_2s60_burst_3_downstream_burstcount),
      .std_2s60_burst_3_downstream_byteenable                     (std_2s60_burst_3_downstream_byteenable),
      .std_2s60_burst_3_downstream_granted_ext_flash_s1           (std_2s60_burst_3_downstream_granted_ext_flash_s1),
      .std_2s60_burst_3_downstream_latency_counter                (std_2s60_burst_3_downstream_latency_counter),
      .std_2s60_burst_3_downstream_qualified_request_ext_flash_s1 (std_2s60_burst_3_downstream_qualified_request_ext_flash_s1),
      .std_2s60_burst_3_downstream_read                           (std_2s60_burst_3_downstream_read),
      .std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1   (std_2s60_burst_3_downstream_read_data_valid_ext_flash_s1),
      .std_2s60_burst_3_downstream_readdata                       (std_2s60_burst_3_downstream_readdata),
      .std_2s60_burst_3_downstream_readdatavalid                  (std_2s60_burst_3_downstream_readdatavalid),
      .std_2s60_burst_3_downstream_requests_ext_flash_s1          (std_2s60_burst_3_downstream_requests_ext_flash_s1),
      .std_2s60_burst_3_downstream_reset_n                        (std_2s60_burst_3_downstream_reset_n),
      .std_2s60_burst_3_downstream_waitrequest                    (std_2s60_burst_3_downstream_waitrequest),
      .std_2s60_burst_3_downstream_write                          (std_2s60_burst_3_downstream_write),
      .std_2s60_burst_3_downstream_writedata                      (std_2s60_burst_3_downstream_writedata)
    );

  std_2s60_burst_3 the_std_2s60_burst_3
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_3_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_3_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_3_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_3_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_3_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_3_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_3_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_3_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_3_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_3_downstream_read),
      .reg_downstream_write            (std_2s60_burst_3_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_3_downstream_writedata),
      .reset_n                         (std_2s60_burst_3_downstream_reset_n),
      .upstream_address                (std_2s60_burst_3_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_3_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_3_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_3_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_3_upstream_address),
      .upstream_read                   (std_2s60_burst_3_upstream_read),
      .upstream_readdata               (std_2s60_burst_3_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_3_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_3_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_3_upstream_write),
      .upstream_writedata              (std_2s60_burst_3_upstream_writedata)
    );

  std_2s60_burst_4_upstream_arbitrator the_std_2s60_burst_4_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_4_upstream                         (cpu_instruction_master_granted_std_2s60_burst_4_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_4_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_4_upstream                        (cpu_instruction_master_requests_std_2s60_burst_4_upstream),
      .d1_std_2s60_burst_4_upstream_end_xfer                                            (d1_std_2s60_burst_4_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_4_upstream_address                                                (std_2s60_burst_4_upstream_address),
      .std_2s60_burst_4_upstream_byteaddress                                            (std_2s60_burst_4_upstream_byteaddress),
      .std_2s60_burst_4_upstream_byteenable                                             (std_2s60_burst_4_upstream_byteenable),
      .std_2s60_burst_4_upstream_debugaccess                                            (std_2s60_burst_4_upstream_debugaccess),
      .std_2s60_burst_4_upstream_read                                                   (std_2s60_burst_4_upstream_read),
      .std_2s60_burst_4_upstream_readdata                                               (std_2s60_burst_4_upstream_readdata),
      .std_2s60_burst_4_upstream_readdata_from_sa                                       (std_2s60_burst_4_upstream_readdata_from_sa),
      .std_2s60_burst_4_upstream_readdatavalid                                          (std_2s60_burst_4_upstream_readdatavalid),
      .std_2s60_burst_4_upstream_waitrequest                                            (std_2s60_burst_4_upstream_waitrequest),
      .std_2s60_burst_4_upstream_waitrequest_from_sa                                    (std_2s60_burst_4_upstream_waitrequest_from_sa),
      .std_2s60_burst_4_upstream_write                                                  (std_2s60_burst_4_upstream_write)
    );

  std_2s60_burst_4_downstream_arbitrator the_std_2s60_burst_4_downstream
    (
      .clk                                                        (clk),
      .d1_ext_ram_bus_avalon_slave_end_xfer                       (d1_ext_ram_bus_avalon_slave_end_xfer),
      .ext_ram_s1_wait_counter_eq_0                               (ext_ram_s1_wait_counter_eq_0),
      .incoming_ext_ram_bus_data                                  (incoming_ext_ram_bus_data),
      .lan91c111_s1_wait_counter_eq_0                             (lan91c111_s1_wait_counter_eq_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_4_downstream_address                        (std_2s60_burst_4_downstream_address),
      .std_2s60_burst_4_downstream_address_to_slave               (std_2s60_burst_4_downstream_address_to_slave),
      .std_2s60_burst_4_downstream_burstcount                     (std_2s60_burst_4_downstream_burstcount),
      .std_2s60_burst_4_downstream_byteenable                     (std_2s60_burst_4_downstream_byteenable),
      .std_2s60_burst_4_downstream_granted_ext_ram_s1             (std_2s60_burst_4_downstream_granted_ext_ram_s1),
      .std_2s60_burst_4_downstream_granted_lan91c111_s1           (std_2s60_burst_4_downstream_granted_lan91c111_s1),
      .std_2s60_burst_4_downstream_latency_counter                (std_2s60_burst_4_downstream_latency_counter),
      .std_2s60_burst_4_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_4_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_4_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_4_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_4_downstream_read                           (std_2s60_burst_4_downstream_read),
      .std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_4_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_4_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_4_downstream_readdata                       (std_2s60_burst_4_downstream_readdata),
      .std_2s60_burst_4_downstream_readdatavalid                  (std_2s60_burst_4_downstream_readdatavalid),
      .std_2s60_burst_4_downstream_requests_ext_ram_s1            (std_2s60_burst_4_downstream_requests_ext_ram_s1),
      .std_2s60_burst_4_downstream_requests_lan91c111_s1          (std_2s60_burst_4_downstream_requests_lan91c111_s1),
      .std_2s60_burst_4_downstream_reset_n                        (std_2s60_burst_4_downstream_reset_n),
      .std_2s60_burst_4_downstream_waitrequest                    (std_2s60_burst_4_downstream_waitrequest),
      .std_2s60_burst_4_downstream_write                          (std_2s60_burst_4_downstream_write),
      .std_2s60_burst_4_downstream_writedata                      (std_2s60_burst_4_downstream_writedata)
    );

  std_2s60_burst_4 the_std_2s60_burst_4
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_4_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_4_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_4_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_4_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_4_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_4_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_4_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_4_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_4_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_4_downstream_read),
      .reg_downstream_write            (std_2s60_burst_4_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_4_downstream_writedata),
      .reset_n                         (std_2s60_burst_4_downstream_reset_n),
      .upstream_address                (std_2s60_burst_4_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_4_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_4_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_4_upstream_address),
      .upstream_read                   (std_2s60_burst_4_upstream_read),
      .upstream_readdata               (std_2s60_burst_4_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_4_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_4_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_4_upstream_write),
      .upstream_writedata              (std_2s60_burst_4_upstream_writedata)
    );

  std_2s60_burst_5_upstream_arbitrator the_std_2s60_burst_5_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_5_upstream                         (cpu_data_master_granted_std_2s60_burst_5_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_5_upstream               (cpu_data_master_qualified_request_std_2s60_burst_5_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_5_upstream                        (cpu_data_master_requests_std_2s60_burst_5_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_5_upstream_end_xfer                                     (d1_std_2s60_burst_5_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_5_upstream_address                                         (std_2s60_burst_5_upstream_address),
      .std_2s60_burst_5_upstream_burstcount                                      (std_2s60_burst_5_upstream_burstcount),
      .std_2s60_burst_5_upstream_byteaddress                                     (std_2s60_burst_5_upstream_byteaddress),
      .std_2s60_burst_5_upstream_byteenable                                      (std_2s60_burst_5_upstream_byteenable),
      .std_2s60_burst_5_upstream_debugaccess                                     (std_2s60_burst_5_upstream_debugaccess),
      .std_2s60_burst_5_upstream_read                                            (std_2s60_burst_5_upstream_read),
      .std_2s60_burst_5_upstream_readdata                                        (std_2s60_burst_5_upstream_readdata),
      .std_2s60_burst_5_upstream_readdata_from_sa                                (std_2s60_burst_5_upstream_readdata_from_sa),
      .std_2s60_burst_5_upstream_readdatavalid                                   (std_2s60_burst_5_upstream_readdatavalid),
      .std_2s60_burst_5_upstream_waitrequest                                     (std_2s60_burst_5_upstream_waitrequest),
      .std_2s60_burst_5_upstream_waitrequest_from_sa                             (std_2s60_burst_5_upstream_waitrequest_from_sa),
      .std_2s60_burst_5_upstream_write                                           (std_2s60_burst_5_upstream_write),
      .std_2s60_burst_5_upstream_writedata                                       (std_2s60_burst_5_upstream_writedata)
    );

  std_2s60_burst_5_downstream_arbitrator the_std_2s60_burst_5_downstream
    (
      .clk                                                        (clk),
      .d1_ext_ram_bus_avalon_slave_end_xfer                       (d1_ext_ram_bus_avalon_slave_end_xfer),
      .ext_ram_s1_wait_counter_eq_0                               (ext_ram_s1_wait_counter_eq_0),
      .incoming_ext_ram_bus_data                                  (incoming_ext_ram_bus_data),
      .lan91c111_s1_wait_counter_eq_0                             (lan91c111_s1_wait_counter_eq_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_5_downstream_address                        (std_2s60_burst_5_downstream_address),
      .std_2s60_burst_5_downstream_address_to_slave               (std_2s60_burst_5_downstream_address_to_slave),
      .std_2s60_burst_5_downstream_burstcount                     (std_2s60_burst_5_downstream_burstcount),
      .std_2s60_burst_5_downstream_byteenable                     (std_2s60_burst_5_downstream_byteenable),
      .std_2s60_burst_5_downstream_granted_ext_ram_s1             (std_2s60_burst_5_downstream_granted_ext_ram_s1),
      .std_2s60_burst_5_downstream_granted_lan91c111_s1           (std_2s60_burst_5_downstream_granted_lan91c111_s1),
      .std_2s60_burst_5_downstream_latency_counter                (std_2s60_burst_5_downstream_latency_counter),
      .std_2s60_burst_5_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_5_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_5_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_5_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_5_downstream_read                           (std_2s60_burst_5_downstream_read),
      .std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_5_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_5_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_5_downstream_readdata                       (std_2s60_burst_5_downstream_readdata),
      .std_2s60_burst_5_downstream_readdatavalid                  (std_2s60_burst_5_downstream_readdatavalid),
      .std_2s60_burst_5_downstream_requests_ext_ram_s1            (std_2s60_burst_5_downstream_requests_ext_ram_s1),
      .std_2s60_burst_5_downstream_requests_lan91c111_s1          (std_2s60_burst_5_downstream_requests_lan91c111_s1),
      .std_2s60_burst_5_downstream_reset_n                        (std_2s60_burst_5_downstream_reset_n),
      .std_2s60_burst_5_downstream_waitrequest                    (std_2s60_burst_5_downstream_waitrequest),
      .std_2s60_burst_5_downstream_write                          (std_2s60_burst_5_downstream_write),
      .std_2s60_burst_5_downstream_writedata                      (std_2s60_burst_5_downstream_writedata)
    );

  std_2s60_burst_5 the_std_2s60_burst_5
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_5_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_5_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_5_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_5_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_5_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_5_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_5_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_5_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_5_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_5_downstream_read),
      .reg_downstream_write            (std_2s60_burst_5_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_5_downstream_writedata),
      .reset_n                         (std_2s60_burst_5_downstream_reset_n),
      .upstream_address                (std_2s60_burst_5_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_5_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_5_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_5_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_5_upstream_address),
      .upstream_read                   (std_2s60_burst_5_upstream_read),
      .upstream_readdata               (std_2s60_burst_5_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_5_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_5_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_5_upstream_write),
      .upstream_writedata              (std_2s60_burst_5_upstream_writedata)
    );

  std_2s60_burst_6_upstream_arbitrator the_std_2s60_burst_6_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_6_upstream                         (cpu_instruction_master_granted_std_2s60_burst_6_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_6_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_6_upstream                        (cpu_instruction_master_requests_std_2s60_burst_6_upstream),
      .d1_std_2s60_burst_6_upstream_end_xfer                                            (d1_std_2s60_burst_6_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_6_upstream_address                                                (std_2s60_burst_6_upstream_address),
      .std_2s60_burst_6_upstream_byteaddress                                            (std_2s60_burst_6_upstream_byteaddress),
      .std_2s60_burst_6_upstream_byteenable                                             (std_2s60_burst_6_upstream_byteenable),
      .std_2s60_burst_6_upstream_debugaccess                                            (std_2s60_burst_6_upstream_debugaccess),
      .std_2s60_burst_6_upstream_read                                                   (std_2s60_burst_6_upstream_read),
      .std_2s60_burst_6_upstream_readdata                                               (std_2s60_burst_6_upstream_readdata),
      .std_2s60_burst_6_upstream_readdata_from_sa                                       (std_2s60_burst_6_upstream_readdata_from_sa),
      .std_2s60_burst_6_upstream_readdatavalid                                          (std_2s60_burst_6_upstream_readdatavalid),
      .std_2s60_burst_6_upstream_waitrequest                                            (std_2s60_burst_6_upstream_waitrequest),
      .std_2s60_burst_6_upstream_waitrequest_from_sa                                    (std_2s60_burst_6_upstream_waitrequest_from_sa),
      .std_2s60_burst_6_upstream_write                                                  (std_2s60_burst_6_upstream_write)
    );

  std_2s60_burst_6_downstream_arbitrator the_std_2s60_burst_6_downstream
    (
      .clk                                                                   (clk),
      .d1_onchip_ram_64_kbytes_s1_end_xfer                                   (d1_onchip_ram_64_kbytes_s1_end_xfer),
      .onchip_ram_64_kbytes_s1_readdata_from_sa                              (onchip_ram_64_kbytes_s1_readdata_from_sa),
      .reset_n                                                               (clk_reset_n),
      .std_2s60_burst_6_downstream_address                                   (std_2s60_burst_6_downstream_address),
      .std_2s60_burst_6_downstream_address_to_slave                          (std_2s60_burst_6_downstream_address_to_slave),
      .std_2s60_burst_6_downstream_burstcount                                (std_2s60_burst_6_downstream_burstcount),
      .std_2s60_burst_6_downstream_byteenable                                (std_2s60_burst_6_downstream_byteenable),
      .std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1           (std_2s60_burst_6_downstream_granted_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_latency_counter                           (std_2s60_burst_6_downstream_latency_counter),
      .std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1 (std_2s60_burst_6_downstream_qualified_request_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_read                                      (std_2s60_burst_6_downstream_read),
      .std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1   (std_2s60_burst_6_downstream_read_data_valid_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_readdata                                  (std_2s60_burst_6_downstream_readdata),
      .std_2s60_burst_6_downstream_readdatavalid                             (std_2s60_burst_6_downstream_readdatavalid),
      .std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1          (std_2s60_burst_6_downstream_requests_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_6_downstream_reset_n                                   (std_2s60_burst_6_downstream_reset_n),
      .std_2s60_burst_6_downstream_waitrequest                               (std_2s60_burst_6_downstream_waitrequest),
      .std_2s60_burst_6_downstream_write                                     (std_2s60_burst_6_downstream_write),
      .std_2s60_burst_6_downstream_writedata                                 (std_2s60_burst_6_downstream_writedata)
    );

  std_2s60_burst_6 the_std_2s60_burst_6
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_6_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_6_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_6_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_6_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_6_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_6_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_6_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_6_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_6_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_6_downstream_read),
      .reg_downstream_write            (std_2s60_burst_6_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_6_downstream_writedata),
      .reset_n                         (std_2s60_burst_6_downstream_reset_n),
      .upstream_address                (std_2s60_burst_6_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_6_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_6_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_6_upstream_address),
      .upstream_read                   (std_2s60_burst_6_upstream_read),
      .upstream_readdata               (std_2s60_burst_6_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_6_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_6_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_6_upstream_write),
      .upstream_writedata              (std_2s60_burst_6_upstream_writedata)
    );

  std_2s60_burst_7_upstream_arbitrator the_std_2s60_burst_7_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_7_upstream                         (cpu_data_master_granted_std_2s60_burst_7_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_7_upstream               (cpu_data_master_qualified_request_std_2s60_burst_7_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_7_upstream                        (cpu_data_master_requests_std_2s60_burst_7_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_7_upstream_end_xfer                                     (d1_std_2s60_burst_7_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_7_upstream_address                                         (std_2s60_burst_7_upstream_address),
      .std_2s60_burst_7_upstream_burstcount                                      (std_2s60_burst_7_upstream_burstcount),
      .std_2s60_burst_7_upstream_byteaddress                                     (std_2s60_burst_7_upstream_byteaddress),
      .std_2s60_burst_7_upstream_byteenable                                      (std_2s60_burst_7_upstream_byteenable),
      .std_2s60_burst_7_upstream_debugaccess                                     (std_2s60_burst_7_upstream_debugaccess),
      .std_2s60_burst_7_upstream_read                                            (std_2s60_burst_7_upstream_read),
      .std_2s60_burst_7_upstream_readdata                                        (std_2s60_burst_7_upstream_readdata),
      .std_2s60_burst_7_upstream_readdata_from_sa                                (std_2s60_burst_7_upstream_readdata_from_sa),
      .std_2s60_burst_7_upstream_readdatavalid                                   (std_2s60_burst_7_upstream_readdatavalid),
      .std_2s60_burst_7_upstream_waitrequest                                     (std_2s60_burst_7_upstream_waitrequest),
      .std_2s60_burst_7_upstream_waitrequest_from_sa                             (std_2s60_burst_7_upstream_waitrequest_from_sa),
      .std_2s60_burst_7_upstream_write                                           (std_2s60_burst_7_upstream_write),
      .std_2s60_burst_7_upstream_writedata                                       (std_2s60_burst_7_upstream_writedata)
    );

  std_2s60_burst_7_downstream_arbitrator the_std_2s60_burst_7_downstream
    (
      .clk                                                                   (clk),
      .d1_onchip_ram_64_kbytes_s1_end_xfer                                   (d1_onchip_ram_64_kbytes_s1_end_xfer),
      .onchip_ram_64_kbytes_s1_readdata_from_sa                              (onchip_ram_64_kbytes_s1_readdata_from_sa),
      .reset_n                                                               (clk_reset_n),
      .std_2s60_burst_7_downstream_address                                   (std_2s60_burst_7_downstream_address),
      .std_2s60_burst_7_downstream_address_to_slave                          (std_2s60_burst_7_downstream_address_to_slave),
      .std_2s60_burst_7_downstream_burstcount                                (std_2s60_burst_7_downstream_burstcount),
      .std_2s60_burst_7_downstream_byteenable                                (std_2s60_burst_7_downstream_byteenable),
      .std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1           (std_2s60_burst_7_downstream_granted_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_latency_counter                           (std_2s60_burst_7_downstream_latency_counter),
      .std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1 (std_2s60_burst_7_downstream_qualified_request_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_read                                      (std_2s60_burst_7_downstream_read),
      .std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1   (std_2s60_burst_7_downstream_read_data_valid_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_readdata                                  (std_2s60_burst_7_downstream_readdata),
      .std_2s60_burst_7_downstream_readdatavalid                             (std_2s60_burst_7_downstream_readdatavalid),
      .std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1          (std_2s60_burst_7_downstream_requests_onchip_ram_64_kbytes_s1),
      .std_2s60_burst_7_downstream_reset_n                                   (std_2s60_burst_7_downstream_reset_n),
      .std_2s60_burst_7_downstream_waitrequest                               (std_2s60_burst_7_downstream_waitrequest),
      .std_2s60_burst_7_downstream_write                                     (std_2s60_burst_7_downstream_write),
      .std_2s60_burst_7_downstream_writedata                                 (std_2s60_burst_7_downstream_writedata)
    );

  std_2s60_burst_7 the_std_2s60_burst_7
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_7_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_7_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_7_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_7_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_7_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_7_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_7_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_7_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_7_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_7_downstream_read),
      .reg_downstream_write            (std_2s60_burst_7_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_7_downstream_writedata),
      .reset_n                         (std_2s60_burst_7_downstream_reset_n),
      .upstream_address                (std_2s60_burst_7_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_7_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_7_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_7_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_7_upstream_address),
      .upstream_read                   (std_2s60_burst_7_upstream_read),
      .upstream_readdata               (std_2s60_burst_7_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_7_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_7_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_7_upstream_write),
      .upstream_writedata              (std_2s60_burst_7_upstream_writedata)
    );

  std_2s60_burst_8_upstream_arbitrator the_std_2s60_burst_8_upstream
    (
      .clk                                                                              (clk),
      .cpu_instruction_master_address_to_slave                                          (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_std_2s60_burst_8_upstream                         (cpu_instruction_master_granted_std_2s60_burst_8_upstream),
      .cpu_instruction_master_latency_counter                                           (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream               (cpu_instruction_master_qualified_request_std_2s60_burst_8_upstream),
      .cpu_instruction_master_read                                                      (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_0_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_15_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register (cpu_instruction_master_read_data_valid_std_2s60_burst_18_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_2_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_4_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_6_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream                 (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream),
      .cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register  (cpu_instruction_master_read_data_valid_std_2s60_burst_8_upstream_shift_register),
      .cpu_instruction_master_requests_std_2s60_burst_8_upstream                        (cpu_instruction_master_requests_std_2s60_burst_8_upstream),
      .d1_std_2s60_burst_8_upstream_end_xfer                                            (d1_std_2s60_burst_8_upstream_end_xfer),
      .reset_n                                                                          (clk_reset_n),
      .std_2s60_burst_8_upstream_address                                                (std_2s60_burst_8_upstream_address),
      .std_2s60_burst_8_upstream_byteaddress                                            (std_2s60_burst_8_upstream_byteaddress),
      .std_2s60_burst_8_upstream_byteenable                                             (std_2s60_burst_8_upstream_byteenable),
      .std_2s60_burst_8_upstream_debugaccess                                            (std_2s60_burst_8_upstream_debugaccess),
      .std_2s60_burst_8_upstream_read                                                   (std_2s60_burst_8_upstream_read),
      .std_2s60_burst_8_upstream_readdata                                               (std_2s60_burst_8_upstream_readdata),
      .std_2s60_burst_8_upstream_readdata_from_sa                                       (std_2s60_burst_8_upstream_readdata_from_sa),
      .std_2s60_burst_8_upstream_readdatavalid                                          (std_2s60_burst_8_upstream_readdatavalid),
      .std_2s60_burst_8_upstream_waitrequest                                            (std_2s60_burst_8_upstream_waitrequest),
      .std_2s60_burst_8_upstream_waitrequest_from_sa                                    (std_2s60_burst_8_upstream_waitrequest_from_sa),
      .std_2s60_burst_8_upstream_write                                                  (std_2s60_burst_8_upstream_write)
    );

  std_2s60_burst_8_downstream_arbitrator the_std_2s60_burst_8_downstream
    (
      .clk                                                        (clk),
      .d1_ext_ram_bus_avalon_slave_end_xfer                       (d1_ext_ram_bus_avalon_slave_end_xfer),
      .ext_ram_s1_wait_counter_eq_0                               (ext_ram_s1_wait_counter_eq_0),
      .incoming_ext_ram_bus_data                                  (incoming_ext_ram_bus_data),
      .lan91c111_s1_wait_counter_eq_0                             (lan91c111_s1_wait_counter_eq_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_8_downstream_address                        (std_2s60_burst_8_downstream_address),
      .std_2s60_burst_8_downstream_address_to_slave               (std_2s60_burst_8_downstream_address_to_slave),
      .std_2s60_burst_8_downstream_burstcount                     (std_2s60_burst_8_downstream_burstcount),
      .std_2s60_burst_8_downstream_byteenable                     (std_2s60_burst_8_downstream_byteenable),
      .std_2s60_burst_8_downstream_granted_ext_ram_s1             (std_2s60_burst_8_downstream_granted_ext_ram_s1),
      .std_2s60_burst_8_downstream_granted_lan91c111_s1           (std_2s60_burst_8_downstream_granted_lan91c111_s1),
      .std_2s60_burst_8_downstream_latency_counter                (std_2s60_burst_8_downstream_latency_counter),
      .std_2s60_burst_8_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_8_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_8_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_8_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_8_downstream_read                           (std_2s60_burst_8_downstream_read),
      .std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_8_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_8_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_8_downstream_readdata                       (std_2s60_burst_8_downstream_readdata),
      .std_2s60_burst_8_downstream_readdatavalid                  (std_2s60_burst_8_downstream_readdatavalid),
      .std_2s60_burst_8_downstream_requests_ext_ram_s1            (std_2s60_burst_8_downstream_requests_ext_ram_s1),
      .std_2s60_burst_8_downstream_requests_lan91c111_s1          (std_2s60_burst_8_downstream_requests_lan91c111_s1),
      .std_2s60_burst_8_downstream_reset_n                        (std_2s60_burst_8_downstream_reset_n),
      .std_2s60_burst_8_downstream_waitrequest                    (std_2s60_burst_8_downstream_waitrequest),
      .std_2s60_burst_8_downstream_write                          (std_2s60_burst_8_downstream_write),
      .std_2s60_burst_8_downstream_writedata                      (std_2s60_burst_8_downstream_writedata)
    );

  std_2s60_burst_8 the_std_2s60_burst_8
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_8_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_8_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_8_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_8_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_8_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_8_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_8_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_8_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_8_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_8_downstream_read),
      .reg_downstream_write            (std_2s60_burst_8_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_8_downstream_writedata),
      .reset_n                         (std_2s60_burst_8_downstream_reset_n),
      .upstream_address                (std_2s60_burst_8_upstream_byteaddress),
      .upstream_byteenable             (std_2s60_burst_8_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_8_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_8_upstream_address),
      .upstream_read                   (std_2s60_burst_8_upstream_read),
      .upstream_readdata               (std_2s60_burst_8_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_8_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_8_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_8_upstream_write),
      .upstream_writedata              (std_2s60_burst_8_upstream_writedata)
    );

  std_2s60_burst_9_upstream_arbitrator the_std_2s60_burst_9_upstream
    (
      .clk                                                                       (clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_std_2s60_burst_9_upstream                         (cpu_data_master_granted_std_2s60_burst_9_upstream),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_std_2s60_burst_9_upstream               (cpu_data_master_qualified_request_std_2s60_burst_9_upstream),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_10_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_11_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_12_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_13_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_14_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_16_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register (cpu_data_master_read_data_valid_std_2s60_burst_17_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_1_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_3_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_5_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_7_upstream_shift_register),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream                 (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream),
      .cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register  (cpu_data_master_read_data_valid_std_2s60_burst_9_upstream_shift_register),
      .cpu_data_master_requests_std_2s60_burst_9_upstream                        (cpu_data_master_requests_std_2s60_burst_9_upstream),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_std_2s60_burst_9_upstream_end_xfer                                     (d1_std_2s60_burst_9_upstream_end_xfer),
      .reset_n                                                                   (clk_reset_n),
      .std_2s60_burst_9_upstream_address                                         (std_2s60_burst_9_upstream_address),
      .std_2s60_burst_9_upstream_burstcount                                      (std_2s60_burst_9_upstream_burstcount),
      .std_2s60_burst_9_upstream_byteaddress                                     (std_2s60_burst_9_upstream_byteaddress),
      .std_2s60_burst_9_upstream_byteenable                                      (std_2s60_burst_9_upstream_byteenable),
      .std_2s60_burst_9_upstream_debugaccess                                     (std_2s60_burst_9_upstream_debugaccess),
      .std_2s60_burst_9_upstream_read                                            (std_2s60_burst_9_upstream_read),
      .std_2s60_burst_9_upstream_readdata                                        (std_2s60_burst_9_upstream_readdata),
      .std_2s60_burst_9_upstream_readdata_from_sa                                (std_2s60_burst_9_upstream_readdata_from_sa),
      .std_2s60_burst_9_upstream_readdatavalid                                   (std_2s60_burst_9_upstream_readdatavalid),
      .std_2s60_burst_9_upstream_waitrequest                                     (std_2s60_burst_9_upstream_waitrequest),
      .std_2s60_burst_9_upstream_waitrequest_from_sa                             (std_2s60_burst_9_upstream_waitrequest_from_sa),
      .std_2s60_burst_9_upstream_write                                           (std_2s60_burst_9_upstream_write),
      .std_2s60_burst_9_upstream_writedata                                       (std_2s60_burst_9_upstream_writedata)
    );

  std_2s60_burst_9_downstream_arbitrator the_std_2s60_burst_9_downstream
    (
      .clk                                                        (clk),
      .d1_ext_ram_bus_avalon_slave_end_xfer                       (d1_ext_ram_bus_avalon_slave_end_xfer),
      .ext_ram_s1_wait_counter_eq_0                               (ext_ram_s1_wait_counter_eq_0),
      .incoming_ext_ram_bus_data                                  (incoming_ext_ram_bus_data),
      .lan91c111_s1_wait_counter_eq_0                             (lan91c111_s1_wait_counter_eq_0),
      .reset_n                                                    (clk_reset_n),
      .std_2s60_burst_9_downstream_address                        (std_2s60_burst_9_downstream_address),
      .std_2s60_burst_9_downstream_address_to_slave               (std_2s60_burst_9_downstream_address_to_slave),
      .std_2s60_burst_9_downstream_burstcount                     (std_2s60_burst_9_downstream_burstcount),
      .std_2s60_burst_9_downstream_byteenable                     (std_2s60_burst_9_downstream_byteenable),
      .std_2s60_burst_9_downstream_granted_ext_ram_s1             (std_2s60_burst_9_downstream_granted_ext_ram_s1),
      .std_2s60_burst_9_downstream_granted_lan91c111_s1           (std_2s60_burst_9_downstream_granted_lan91c111_s1),
      .std_2s60_burst_9_downstream_latency_counter                (std_2s60_burst_9_downstream_latency_counter),
      .std_2s60_burst_9_downstream_qualified_request_ext_ram_s1   (std_2s60_burst_9_downstream_qualified_request_ext_ram_s1),
      .std_2s60_burst_9_downstream_qualified_request_lan91c111_s1 (std_2s60_burst_9_downstream_qualified_request_lan91c111_s1),
      .std_2s60_burst_9_downstream_read                           (std_2s60_burst_9_downstream_read),
      .std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1     (std_2s60_burst_9_downstream_read_data_valid_ext_ram_s1),
      .std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1   (std_2s60_burst_9_downstream_read_data_valid_lan91c111_s1),
      .std_2s60_burst_9_downstream_readdata                       (std_2s60_burst_9_downstream_readdata),
      .std_2s60_burst_9_downstream_readdatavalid                  (std_2s60_burst_9_downstream_readdatavalid),
      .std_2s60_burst_9_downstream_requests_ext_ram_s1            (std_2s60_burst_9_downstream_requests_ext_ram_s1),
      .std_2s60_burst_9_downstream_requests_lan91c111_s1          (std_2s60_burst_9_downstream_requests_lan91c111_s1),
      .std_2s60_burst_9_downstream_reset_n                        (std_2s60_burst_9_downstream_reset_n),
      .std_2s60_burst_9_downstream_waitrequest                    (std_2s60_burst_9_downstream_waitrequest),
      .std_2s60_burst_9_downstream_write                          (std_2s60_burst_9_downstream_write),
      .std_2s60_burst_9_downstream_writedata                      (std_2s60_burst_9_downstream_writedata)
    );

  std_2s60_burst_9 the_std_2s60_burst_9
    (
      .clk                             (clk),
      .downstream_readdata             (std_2s60_burst_9_downstream_readdata),
      .downstream_readdatavalid        (std_2s60_burst_9_downstream_readdatavalid),
      .downstream_waitrequest          (std_2s60_burst_9_downstream_waitrequest),
      .reg_downstream_address          (std_2s60_burst_9_downstream_address),
      .reg_downstream_arbitrationshare (std_2s60_burst_9_downstream_arbitrationshare),
      .reg_downstream_burstcount       (std_2s60_burst_9_downstream_burstcount),
      .reg_downstream_byteenable       (std_2s60_burst_9_downstream_byteenable),
      .reg_downstream_debugaccess      (std_2s60_burst_9_downstream_debugaccess),
      .reg_downstream_nativeaddress    (std_2s60_burst_9_downstream_nativeaddress),
      .reg_downstream_read             (std_2s60_burst_9_downstream_read),
      .reg_downstream_write            (std_2s60_burst_9_downstream_write),
      .reg_downstream_writedata        (std_2s60_burst_9_downstream_writedata),
      .reset_n                         (std_2s60_burst_9_downstream_reset_n),
      .upstream_address                (std_2s60_burst_9_upstream_byteaddress),
      .upstream_burstcount             (std_2s60_burst_9_upstream_burstcount),
      .upstream_byteenable             (std_2s60_burst_9_upstream_byteenable),
      .upstream_debugaccess            (std_2s60_burst_9_upstream_debugaccess),
      .upstream_nativeaddress          (std_2s60_burst_9_upstream_address),
      .upstream_read                   (std_2s60_burst_9_upstream_read),
      .upstream_readdata               (std_2s60_burst_9_upstream_readdata),
      .upstream_readdatavalid          (std_2s60_burst_9_upstream_readdatavalid),
      .upstream_waitrequest            (std_2s60_burst_9_upstream_waitrequest),
      .upstream_write                  (std_2s60_burst_9_upstream_write),
      .upstream_writedata              (std_2s60_burst_9_upstream_writedata)
    );

  sys_clk_timer_s1_arbitrator the_sys_clk_timer_s1
    (
      .clk                                                             (clk),
      .d1_sys_clk_timer_s1_end_xfer                                    (d1_sys_clk_timer_s1_end_xfer),
      .reset_n                                                         (clk_reset_n),
      .std_2s60_burst_10_downstream_address_to_slave                   (std_2s60_burst_10_downstream_address_to_slave),
      .std_2s60_burst_10_downstream_arbitrationshare                   (std_2s60_burst_10_downstream_arbitrationshare),
      .std_2s60_burst_10_downstream_burstcount                         (std_2s60_burst_10_downstream_burstcount),
      .std_2s60_burst_10_downstream_granted_sys_clk_timer_s1           (std_2s60_burst_10_downstream_granted_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_latency_counter                    (std_2s60_burst_10_downstream_latency_counter),
      .std_2s60_burst_10_downstream_nativeaddress                      (std_2s60_burst_10_downstream_nativeaddress),
      .std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1 (std_2s60_burst_10_downstream_qualified_request_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_read                               (std_2s60_burst_10_downstream_read),
      .std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1   (std_2s60_burst_10_downstream_read_data_valid_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_requests_sys_clk_timer_s1          (std_2s60_burst_10_downstream_requests_sys_clk_timer_s1),
      .std_2s60_burst_10_downstream_write                              (std_2s60_burst_10_downstream_write),
      .std_2s60_burst_10_downstream_writedata                          (std_2s60_burst_10_downstream_writedata),
      .sys_clk_timer_s1_address                                        (sys_clk_timer_s1_address),
      .sys_clk_timer_s1_chipselect                                     (sys_clk_timer_s1_chipselect),
      .sys_clk_timer_s1_irq                                            (sys_clk_timer_s1_irq),
      .sys_clk_timer_s1_irq_from_sa                                    (sys_clk_timer_s1_irq_from_sa),
      .sys_clk_timer_s1_readdata                                       (sys_clk_timer_s1_readdata),
      .sys_clk_timer_s1_readdata_from_sa                               (sys_clk_timer_s1_readdata_from_sa),
      .sys_clk_timer_s1_reset_n                                        (sys_clk_timer_s1_reset_n),
      .sys_clk_timer_s1_write_n                                        (sys_clk_timer_s1_write_n),
      .sys_clk_timer_s1_writedata                                      (sys_clk_timer_s1_writedata)
    );

  sys_clk_timer the_sys_clk_timer
    (
      .address    (sys_clk_timer_s1_address),
      .chipselect (sys_clk_timer_s1_chipselect),
      .clk        (clk),
      .irq        (sys_clk_timer_s1_irq),
      .readdata   (sys_clk_timer_s1_readdata),
      .reset_n    (sys_clk_timer_s1_reset_n),
      .write_n    (sys_clk_timer_s1_write_n),
      .writedata  (sys_clk_timer_s1_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                                (clk),
      .d1_sysid_control_slave_end_xfer                                    (d1_sysid_control_slave_end_xfer),
      .reset_n                                                            (clk_reset_n),
      .std_2s60_burst_14_downstream_address_to_slave                      (std_2s60_burst_14_downstream_address_to_slave),
      .std_2s60_burst_14_downstream_arbitrationshare                      (std_2s60_burst_14_downstream_arbitrationshare),
      .std_2s60_burst_14_downstream_burstcount                            (std_2s60_burst_14_downstream_burstcount),
      .std_2s60_burst_14_downstream_granted_sysid_control_slave           (std_2s60_burst_14_downstream_granted_sysid_control_slave),
      .std_2s60_burst_14_downstream_latency_counter                       (std_2s60_burst_14_downstream_latency_counter),
      .std_2s60_burst_14_downstream_nativeaddress                         (std_2s60_burst_14_downstream_nativeaddress),
      .std_2s60_burst_14_downstream_qualified_request_sysid_control_slave (std_2s60_burst_14_downstream_qualified_request_sysid_control_slave),
      .std_2s60_burst_14_downstream_read                                  (std_2s60_burst_14_downstream_read),
      .std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave   (std_2s60_burst_14_downstream_read_data_valid_sysid_control_slave),
      .std_2s60_burst_14_downstream_requests_sysid_control_slave          (std_2s60_burst_14_downstream_requests_sysid_control_slave),
      .std_2s60_burst_14_downstream_write                                 (std_2s60_burst_14_downstream_write),
      .sysid_control_slave_address                                        (sysid_control_slave_address),
      .sysid_control_slave_readdata                                       (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                               (sysid_control_slave_readdata_from_sa)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .readdata (sysid_control_slave_readdata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  std_2s60_reset_clk_domain_synch_module std_2s60_reset_clk_domain_synch
    (
      .clk      (clk),
      .data_in  (1'b1),
      .data_out (clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa);

  //std_2s60_burst_0_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_0_upstream_writedata = 0;

  //std_2s60_burst_15_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_15_upstream_writedata = 0;

  //std_2s60_burst_18_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_18_upstream_writedata = 0;

  //std_2s60_burst_2_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_2_upstream_writedata = 0;

  //std_2s60_burst_4_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_4_upstream_writedata = 0;

  //std_2s60_burst_6_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_6_upstream_writedata = 0;

  //std_2s60_burst_8_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign std_2s60_burst_8_upstream_writedata = 0;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane0_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [16777215: 0];
  wire    [  7: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      if (1)
          read_address <= rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      if (1)
//          read_address <= rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash (
                   // inputs:
                    address,
                    read_n,
                    select_n,
                    write_n,

                   // outputs:
                    data
                 )
;

  inout   [  7: 0] data;
  input   [ 23: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [  7: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_flash_lane0, which is an e_ram
  ext_flash_lane0_module ext_flash_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? q_0: {8{1'bz}};

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_lane0_module (
                              // inputs:
                               data,
                               rdaddress,
                               rdclken,
                               wraddress,
                               wrclock,
                               wren,

                              // outputs:
                               q
                            )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      if (1)
          read_address <= rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ram_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      if (1)
//          read_address <= rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ram_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_lane1_module (
                              // inputs:
                               data,
                               rdaddress,
                               rdclken,
                               wraddress,
                               wrclock,
                               wren,

                              // outputs:
                               q
                            )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      if (1)
          read_address <= rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ram_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      if (1)
//          read_address <= rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ram_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_lane2_module (
                              // inputs:
                               data,
                               rdaddress,
                               rdclken,
                               wraddress,
                               wrclock,
                               wren,

                              // outputs:
                               q
                            )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      if (1)
          read_address <= rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ram_lane2.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      if (1)
//          read_address <= rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ram_lane2.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram_lane3_module (
                              // inputs:
                               data,
                               rdaddress,
                               rdclken,
                               wraddress,
                               wrclock,
                               wren,

                              // outputs:
                               q
                            )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      if (1)
          read_address <= rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ram_lane3.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      if (1)
//          read_address <= rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ram_lane3.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ram (
                 // inputs:
                  address,
                  be_n,
                  read_n,
                  select_n,
                  write_n,

                 // outputs:
                  data
               )
;

  inout   [ 31: 0] data;
  input   [ 17: 0] address;
  input   [  3: 0] be_n;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 31: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [  7: 0] data_2;
  wire    [  7: 0] data_3;
  wire    [ 31: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  wire    [  7: 0] q_2;
  wire    [  7: 0] q_3;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_ram_lane0, which is an e_ram
  ext_ram_lane0_module ext_ram_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n & ~be_n[0])
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_ram_lane1, which is an e_ram
  ext_ram_lane1_module ext_ram_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n & ~be_n[1])
    );

  assign data_2 = logic_vector_gasket[23 : 16];
  //ext_ram_lane2, which is an e_ram
  ext_ram_lane2_module ext_ram_lane2
    (
      .data      (data_2),
      .q         (q_2),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n & ~be_n[2])
    );

  assign data_3 = logic_vector_gasket[31 : 24];
  //ext_ram_lane3, which is an e_ram
  ext_ram_lane3_module ext_ram_lane3
    (
      .data      (data_3),
      .q         (q_3),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n & ~be_n[3])
    );

  assign data = (~select_n & ~read_n)? {q_3,
    q_2,
    q_1,
    q_0}: {32{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "c:/altera/quartus80/quartus/eda/sim_lib/altera_mf.v"
`include "c:/altera/quartus80/quartus/eda/sim_lib/220model.v"
`include "c:/altera/quartus80/quartus/eda/sim_lib/sgate.v"
`include "ad_buf.v"
`include "adBUF.v"
`include "std_2s60_burst_17.v"
`include "sdram.v"
`include "sdram_test_component.v"
`include "sysid.v"
`include "high_res_timer.v"
`include "std_2s60_burst_18.v"
`include "std_2s60_burst_13.v"
`include "std_2s60_burst_9.v"
`include "jtag_uart.v"
`include "std_2s60_burst_16.v"
`include "reconfig_request_pio.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "onchip_ram_64_kbytes.v"
`include "std_2s60_burst_4.v"
`include "std_2s60_burst_12.v"
`include "std_2s60_burst_5.v"
`include "std_2s60_burst_3.v"
`include "std_2s60_burst_7.v"
`include "std_2s60_burst_1.v"
`include "std_2s60_burst_0.v"
`include "std_2s60_burst_2.v"
`include "std_2s60_burst_10.v"
`include "sys_clk_timer.v"
`include "std_2s60_burst_11.v"
`include "std_2s60_burst_14.v"
`include "std_2s60_burst_6.v"
`include "std_2s60_burst_8.v"
`include "std_2s60_burst_15.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire    [ 11: 0] a2dc_to_the_ad_buf;
  wire             adclk_to_the_ad_buf;
  wire    [  3: 0] be_n_to_the_ext_ram;
  wire             bidir_port_to_and_from_the_reconfig_request_pio;
  reg              clk;
  wire    [ 23: 0] ext_flash_bus_address;
  wire    [  7: 0] ext_flash_bus_data;
  wire             ext_flash_bus_readn;
  wire    [ 19: 0] ext_ram_bus_address;
  wire    [  3: 0] ext_ram_bus_byteenablen;
  wire    [ 31: 0] ext_ram_bus_data;
  wire             ior_n_to_the_lan91c111;
  wire             iow_n_to_the_lan91c111;
  wire             irq_from_the_lan91c111;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             read_n_to_the_ext_ram;
  reg              reset_n;
  wire             reset_to_the_lan91c111;
  wire             select_n_to_the_ext_flash;
  wire             select_n_to_the_ext_ram;
  wire    [ 10: 0] std_2s60_burst_0_downstream_nativeaddress;
  wire    [ 31: 0] std_2s60_burst_0_upstream_writedata;
  wire             std_2s60_burst_10_downstream_debugaccess;
  wire             std_2s60_burst_11_downstream_debugaccess;
  wire             std_2s60_burst_12_downstream_debugaccess;
  wire             std_2s60_burst_13_downstream_debugaccess;
  wire             std_2s60_burst_14_downstream_debugaccess;
  wire             std_2s60_burst_15_downstream_debugaccess;
  wire    [ 23: 0] std_2s60_burst_15_downstream_nativeaddress;
  wire    [ 31: 0] std_2s60_burst_15_upstream_writedata;
  wire             std_2s60_burst_16_downstream_debugaccess;
  wire    [ 23: 0] std_2s60_burst_16_downstream_nativeaddress;
  wire             std_2s60_burst_17_downstream_debugaccess;
  wire    [ 13: 0] std_2s60_burst_17_downstream_nativeaddress;
  wire             std_2s60_burst_18_downstream_debugaccess;
  wire    [ 13: 0] std_2s60_burst_18_downstream_nativeaddress;
  wire    [ 31: 0] std_2s60_burst_18_upstream_writedata;
  wire    [ 10: 0] std_2s60_burst_1_downstream_nativeaddress;
  wire             std_2s60_burst_2_downstream_debugaccess;
  wire    [ 23: 0] std_2s60_burst_2_downstream_nativeaddress;
  wire    [  7: 0] std_2s60_burst_2_upstream_writedata;
  wire             std_2s60_burst_3_downstream_debugaccess;
  wire    [ 23: 0] std_2s60_burst_3_downstream_nativeaddress;
  wire             std_2s60_burst_4_downstream_debugaccess;
  wire    [ 31: 0] std_2s60_burst_4_upstream_writedata;
  wire             std_2s60_burst_5_downstream_debugaccess;
  wire             std_2s60_burst_6_downstream_debugaccess;
  wire    [ 15: 0] std_2s60_burst_6_downstream_nativeaddress;
  wire    [ 31: 0] std_2s60_burst_6_upstream_writedata;
  wire             std_2s60_burst_7_downstream_debugaccess;
  wire    [ 15: 0] std_2s60_burst_7_downstream_nativeaddress;
  wire             std_2s60_burst_8_downstream_debugaccess;
  wire    [ 31: 0] std_2s60_burst_8_upstream_writedata;
  wire             std_2s60_burst_9_downstream_debugaccess;
  wire             wrclk_to_the_ad_buf;
  wire             write_n_to_the_ext_flash;
  wire             write_n_to_the_ext_ram;
  wire    [ 11: 0] zs_addr_from_the_sdram;
  wire    [  1: 0] zs_ba_from_the_sdram;
  wire             zs_cas_n_from_the_sdram;
  wire             zs_cke_from_the_sdram;
  wire             zs_cs_n_from_the_sdram;
  wire    [ 31: 0] zs_dq_to_and_from_the_sdram;
  wire    [  3: 0] zs_dqm_from_the_sdram;
  wire             zs_ras_n_from_the_sdram;
  wire             zs_we_n_from_the_sdram;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  std_2s60 DUT
    (
      .a2dc_to_the_ad_buf                              (a2dc_to_the_ad_buf),
      .adclk_to_the_ad_buf                             (adclk_to_the_ad_buf),
      .be_n_to_the_ext_ram                             (be_n_to_the_ext_ram),
      .bidir_port_to_and_from_the_reconfig_request_pio (bidir_port_to_and_from_the_reconfig_request_pio),
      .clk                                             (clk),
      .ext_flash_bus_address                           (ext_flash_bus_address),
      .ext_flash_bus_data                              (ext_flash_bus_data),
      .ext_flash_bus_readn                             (ext_flash_bus_readn),
      .ext_ram_bus_address                             (ext_ram_bus_address),
      .ext_ram_bus_byteenablen                         (ext_ram_bus_byteenablen),
      .ext_ram_bus_data                                (ext_ram_bus_data),
      .ior_n_to_the_lan91c111                          (ior_n_to_the_lan91c111),
      .iow_n_to_the_lan91c111                          (iow_n_to_the_lan91c111),
      .irq_from_the_lan91c111                          (irq_from_the_lan91c111),
      .read_n_to_the_ext_ram                           (read_n_to_the_ext_ram),
      .reset_n                                         (reset_n),
      .reset_to_the_lan91c111                          (reset_to_the_lan91c111),
      .select_n_to_the_ext_flash                       (select_n_to_the_ext_flash),
      .select_n_to_the_ext_ram                         (select_n_to_the_ext_ram),
      .wrclk_to_the_ad_buf                             (wrclk_to_the_ad_buf),
      .write_n_to_the_ext_flash                        (write_n_to_the_ext_flash),
      .write_n_to_the_ext_ram                          (write_n_to_the_ext_ram),
      .zs_addr_from_the_sdram                          (zs_addr_from_the_sdram),
      .zs_ba_from_the_sdram                            (zs_ba_from_the_sdram),
      .zs_cas_n_from_the_sdram                         (zs_cas_n_from_the_sdram),
      .zs_cke_from_the_sdram                           (zs_cke_from_the_sdram),
      .zs_cs_n_from_the_sdram                          (zs_cs_n_from_the_sdram),
      .zs_dq_to_and_from_the_sdram                     (zs_dq_to_and_from_the_sdram),
      .zs_dqm_from_the_sdram                           (zs_dqm_from_the_sdram),
      .zs_ras_n_from_the_sdram                         (zs_ras_n_from_the_sdram),
      .zs_we_n_from_the_sdram                          (zs_we_n_from_the_sdram)
    );

  ext_flash the_ext_flash
    (
      .address  (ext_flash_bus_address),
      .data     (ext_flash_bus_data),
      .read_n   (ext_flash_bus_readn),
      .select_n (select_n_to_the_ext_flash),
      .write_n  (write_n_to_the_ext_flash)
    );

  ext_ram the_ext_ram
    (
      .address  (ext_ram_bus_address[19 : 2]),
      .be_n     (be_n_to_the_ext_ram),
      .data     (ext_ram_bus_data),
      .read_n   (read_n_to_the_ext_ram),
      .select_n (select_n_to_the_ext_ram),
      .write_n  (write_n_to_the_ext_ram)
    );

  //default value specified in MODULE lan91c111 ptf port section
  assign irq_from_the_lan91c111 = 0;

  sdram_test_component the_sdram_test_component
    (
      .clk      (clk),
      .zs_addr  (zs_addr_from_the_sdram),
      .zs_ba    (zs_ba_from_the_sdram),
      .zs_cas_n (zs_cas_n_from_the_sdram),
      .zs_cke   (zs_cke_from_the_sdram),
      .zs_cs_n  (zs_cs_n_from_the_sdram),
      .zs_dq    (zs_dq_to_and_from_the_sdram),
      .zs_dqm   (zs_dqm_from_the_sdram),
      .zs_ras_n (zs_ras_n_from_the_sdram),
      .zs_we_n  (zs_we_n_from_the_sdram)
    );

  initial
    clk = 1'b0;
  always
    #3 clk <= ~clk;
  
  initial 
    begin
      reset_n <= 0;
      #65 reset_n <= 1;
    end

endmodule


//synthesis translate_on