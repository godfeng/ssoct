��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��W N��|C��#�N' ���x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`h��>��ׯ�=>)m��U���T���딣0&_���X0���2|	p��rw@	@us���XH����U��h�`.yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|+��@-�-'P�e`b�T=폳�H?o7\F���r��RL�a)�ƞ��U<N	:.���n��{�'����������7C��Hq-/��@�]\���<��9�`J�=�OLl??�L��y�����c��(r���U��óL=��+/��aG�k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Qe�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3"C��dKBE	�\�Z�م�L�Xڈ*-��]���P��`�.�D���J7"~����d6�Pr"?D2BC��5��Yk"1/���%	v3"C��dKBE�磋��w.V&��B֥�(����5���.�^�9��ǘ^�?�;��XC�,�-fce��,\ަ�It�k\,آ(&l�����W����\�v�T?�7G|`h�' L� U��֜��3�LH$��^��{�OF8%v@����fct�:��RE��ʐx�?ێ
7�\Z9�	��%т��!o.sG[�� �tS���}�#�ڊ<?@��[	J��;ι��QG�����U��7�ܥ��2�\Z�ؿH�j�\|Z��0[����	��N�Ae�#�̲�2�!������5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�^�9.�JQ�����5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�eן�-�Q�Z�pMݦ�l��-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0Tu�q�.:�TD��m�jp=�#{��p�{&l����_::���4�ˈ<�I7��-5��6��	���`y������_۾�k�����5	��]�!����M[��Ǣw�)��O�ҋX����>��l%i�-�M�g������{l�f|�ό���.���|��p��h�d �'���Xw�E�i�m}6*�3���f�]�!���D��L#�6�ǌ�lA�1�:�Ω�"��ұ��:�͟�C���F�N~Y��C�Y�)��NË�����8��z{��E�EYZ/�矘��-n��I�?g�f?2)��ׯ�=>̷�8MS�K�E�\��Y �*��H�q���r�x�\�F���ANʂ�g��U-�e�:`�0&l����P2�$:��ι�����/�X�>���
_�n�@/%{�;���;�L���9o��+hi�?O��K�����=ў@'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,D�=P��[W���D��gl�L��M�,���	N^�U���������GZ>.�0�CyW�f�tR�wX�����/��&��4��)@�<[n^/��u�h����ç;-;*�7��X~J�=��n(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���hY����r��C
'~*��#��ꢗ/}����g�ξ������ei�7#�)z� ��4��)�����
�CӞDOɃ&��BM7�k��9�/��q�&�>��왩�2��� �� Ϳ�$��0z�cUL�n����4���á�~O�"j���b7|#9���b!��u����m�#Y"z�a<�Y�{'%s���'����F�r�f�t��6��	���`y����@����gG�[bGf���;F5@0�Z鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀ�T:���V����/��d�٣��c�A�L'��!�a��5�%]���a(􆿳���2����.��DP֞ �(nyfW��􇃬Tk��A3�(N��㎏qló�Q���l�,�Aٺ�Ha(􆿳���2����.���N$ve����􇃬Tk��A3�(N��㎏qló�Q���l��U����T�\ ��i3�|)sՀ�T:���V�V[�b2�k�:A�	S�r��AR1<I�0�f�#/��=��K���ձ�Z��8���/��O���O��ْ5
�8��S��?�F��SO�P��P����&��B�"p�l~V��o5]��lO ܅d�� л�E��QvfZ!4Я\�rƛ�}���1�)�c��!�`�(i3�E����F�Z�>)�ώ�~+�ݗ����>[H��_0Vձ!�`�(i3,ԯ���gn��Ab�%^��}Dq�f����gRI/)�ak�m6�E����F�Z�>)�����˟y���!s�;�Rn\�_c����L�{���D	��U�l>o��|��P�^/�h���/�dSƏw0���wN��0]fH��>d]=]A��O�T=�4e=��-Y�VN�=�ԕd�tuшb��jߺ��0�5tU���+�J��U<o^.K�}/��<Ӭ��|#HK��@=���b��0�5tUзq8�Ј)w�<�_N`E�cvR+��}Dq�f���R��V���X�&�E����F���8�TP��@E�`�8���&��Ŷ;���I�PD�na"�,�>E��4];ˍH����TI��Ԫ,щ�"��<H��(����O�c����L�{jݭ�F���p� o��]��hy�/B/���^!�������>�s�/���U<o^.K�}qW8+����8���&�qr�^*4y-X��;^�8�1-i4];ˍH��E�(��n6�Ѯ� л�U��v��;fZ!4Я\�rƛ�}��k�-i�9~�!�`�(i3!�`�(i3,ԯ���gn��Ab�%^��}Dq�f��N�v�1��B�r��!�`�(i3,ԯ���gn��Ab�%^��}Dq�f����gRI/,�Xʚ@h!�`�(i3,ԯ���gn�J����� ��}Dq�f�{p�R�I8$vVqYY!�`�(i3���D	��U�l>o��|���JLm|��������A?Љ'�-{<qH�~�!�`�(i37�ܥ��2���kܪ���*�LNm�d�tu���ād�,��x��B5�!�`�(i3x�]�V����:L���2*Q=F��:УWKŃS:H��+܆"BT�(���B�r��зq8�Ј)w�<�_N`E�cvR+��}Dq�f�{p�R�I8��a�=L!�`�(i3���D	��U�l>o��|���bǬ�='�u�uX]�Rn\�_�B�r��"�,�>E��4];ˍH��\B�����g�q~[{Q��`�)J*;�p�aٓ�v1a{J�*�8#�������8�TPm=_g}b��t�֚S��~r�S\w���!�`�(i3зq8�Ј)w�<�_N��M��+?���C&���t� ��Oz!�
�W@!�`�(i3���+�J��U<o^.K�}/��<Ӭ�/�"����J^L��z!�
�W@!�`�(i37�ܥ��2�`e7��9��×�>��|�\m���X����,�Xʚ@h�E����F���8�TP��@E�`�8���&��Ŷ;��z!�
�W@!�`�(i3=]A��O�T=�4e=��-Y�VN�=��7p�J��PWV����ftj5 8��!�`�(i3jݭ�F���p� o��]��hy�/B/���^!�������>,�Xʚ@hx�]�V���t���CՐ3��F<Y��j3��� Q�N��*���������c�] S�4];ˍH��E�(��<���A�� ;�Ӆ�&�`�����k@|�%5'��E����F���8�TP��]&�Hž_�FȘ�i��Nj�,�F�v��@���z\�m���Iϕ������z_۬=�!�`�(i3"�,�>E��4];ˍH�C#��N;F��D]�+�~���{/��I(�c?Hh�`K]!�`�(i3!�`�(i3!�`�(i3jݭ�F���,Y�y^:�3�y��j��k��V��e�LtW��e���d�tAAI�O����07�ܥ��2�k��`����VU��d�˰8���&�-�_��>H��n�-�!�`�(i3!�`�(i3���+�J��U<o^.K�}��HwL�X�|#HK��fu��n�!�`�(i3!�`�(i3!�`�(i3���D	��U�l>o��|���z>�n�S�|#HK��fu��n���H�1�� !�`�(i3!�`�(i3���D	��U�l>o��|���z>�n�S���*y}e��?=�2����o��!�`�(i3!�`�(i3,ԯ���gn�J����� ��}Dq�f���R~�e��ד*�h��F�v�C!�`�(i3=]A��O�T=�4e=��-������yM�8���&�9��^K��[N���b�����sd�!�`�(i3���+�J��U<o^.K�},ufOX�mCž_�FȤo�f�Ԝ��MU�@!~�X����Ѵ���X:��+�
H��m��E4];ˍH��1l��m�ئ��b�􏮚ǖ�!�����T"*�M��d��p∺V��܅���9��ȓM�Me����OA�,s>w��Bw�B�"p�l~/�"���꤭%�3��{�o��C!T*p�VU��J!�`�(i3!�`�(i3!�`�(i3"�,�>E���� &N��nF�d����
F�`�����1݁mP2<WV��
i�c�r�N>�X�5G�7Ê7�E�4'���Xw!�`�(i3!�`�(i3!�`�(i3!�`�(i3)��� ��1����_<X����"�����q��l0+���yn�����門�ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%j!bM�9�&?�>�M�O�IQ���}t�{#	�x�u��߹c���o��C!T*Y�{'%s��F���u@����]�7�v�ԯ��Nb-�h�dN�<@Iv�,.9������:5A��p��1���P�Ivu.rg�q��l0q�\E��0���門�ҋX������S8�=	���/|2��#�	�T�\ ���KD��}[e��0�U�S{����<�6�Q=�qő��{XҹvXI)�vNd�)i�'�al��p�@��O���Z鎬�������(���pu�˂�tj{%��ߛ�8���/���}Dq�f�F�d����k�2��J>eR�<�V�Zt%��m&<�,0 ���Ţ�{l�f|��rs�i���YN���o#�_T��,0=]^	�&Z�n��[��{_8�Y���˂lq�㜯}Dq�f�F�d����4�������eR�<�V�ȓM�Me��aL�!��t�j�!󊾵�e�;Pq]g\ ���ǋҠ7�	�ߥ�H�^ /m�6���<�6�Q=���Ң�Q<�6�Q=	I%Mq��`Ҧ�׶!z1��,,ҹ�$�OD��G͘��P�!а��K��k-J����:M���FM�`;$�l���1��in�uM������A��[B�)�b!F��9�����Ïb�}������c�.D�#�ҒIs{�>Y��}�:_�_5:��(�I>�IP�b������:�kR�$fOyQ���؟�-�X��_��n��&�P��00�Ͷ\��[��=<�6�Q=�w�3����f
�@"��g�����Mgs�4�H�O��	�� ��Fw"�Ş|H��S��q<� �77AƐ^�8�s�٩�삢^��)('���Xw�����U���=����t�kD��*�ҋX����L$�����/���%��Y�i`YS����O0�P2<WV�����F�eO�V2y/��S:�cN���dt�{�Yi`YS����6+W��!�`�(i3!�`�(i3<�6�Q=�U�"���M]�B��5.��$�]��tK�"8���ɮ�� л�B)vظ�u�!�`�(i3!�`�(i3���y��lD�U&"���+c��k��Vj����C$��*V�ֆ�\��[��=��hy�xl��B �i<��z��}�<ͧ�:|�"��ӌ�r,�ttT𔛨Z��ΣS�)37J*u�,�JL���*��c�d}];�SSyZr@u!�0�"� ��w� 9_�똣w�ٽv�yq�`0�|(O��"��"�T�>�#�ҒIs{�D������:_�_5:��(�I>�IP�b�����LQo����������0��]㯟�Ķ��d����;���!�v{:��h�k-J����:M���FM�`;$�l���1��in���� zԻ�弳$_N� ���ui�X\�̈́nlH�I<�6�Q=���x��<�6�Q=	I%Mq��`Ҧ�׶!z1��,���F��qJ�?�̃�*�`��n�E�T����X�=���P�;�ȓM�Me���T��G���X��4tΘIy����ߗ��L1�%TԞ}�{J��n��&�P��k<kbm�t�vc;?N�ʡV�l�竷b��"&�=��(��Z鎬����Ĺ#{����}Dq�f���#:�LH�ҋX����L$�����/�����z|�\m���SLq�N���@��O���Z鎬����Ĺ#{����}Dq�f��5Nleo��ݑ���<��z��}�<ͧ�:|�>d�g�K��I(�c@� ��<��z��}�0z�cUL9kX����_G��?g��ORuD,0=]^	�&Z�n��[��{_8�Y���˂lq�㜯}Dq�f�F�d������~�~�8�1P��#K�SM0.�>k0��0ǽi�*��]�!��	Ǹ�y85��q幊s�?����H�c�B���)�g��U-�ee�@Rv����my$�N��;� ��b�� л�d�q=N$,����hQ���}VA�ڦ�c4�RP�m��q��ˑ��N��k�I#�\(z:�ĭ3S��n��@IE�U����S8�=	���/lg������T�\ �́��Wl� -��J�x"GeY𶣂���S.��TD���rs�i���YN���j[��v2ba(􆿳����r
��qő��{r��  <�!�d�<8�c{}�x���� ��6%j_�z����ҧ���I"�Tv{��lw	>F����D�(%�����Ε3��"%���ۂ�3U�?��)�Rݛ��%�5��lW0۳�*ȑs;��|B����k2��� �����!�`�(i3^�R���c+��;�����$�`V1��eX�:&���!�`�(i3!�`�(i3�gKh�ߕ�ő̓Vo\Ӽ�gy�A�Q�#<4^�?���4�蔖9�Ni�v��Q�P���r�<Uee�,�Aٺ�H���H�V�7�}�!����(����
W�Q�x�ӑ��]�~]'\gWg�i4�\3������+�^n=\f�5>���j����v�۲=�k2!�`�(i3�璓�c�������t �[l;M?��y�!�`�(i32W���R0��h޻_KEP��v{��lw	��f��O���k�җ�w!�`�(i3�5ߧE4�퉅�%>�rG߸��S�ȌM�>Fr���X�ǎs�Ӑg�(O՘�O�q�:뺾�7Z������<�6�o8:4ڎ�\��q�O.C��ݚ�Н�ϝ�j
������h��`�����y_�mS8<�n�ݚ�Н�{k�h�+?��	��٨0�����NW���y�N���At��T��Qm�5���J>n���e�S�[2��� ��y���!�`�(i3"<�GU8o_�mS8<�n�ݚ�Н�,��G��z��At��T��Qm�K�A[}��!�`�(i3�%@��w��7��B1"�G!�`�(i3!�`�(i3����P`��]5�d�4䋭�`Z���Y��(�R��#H+�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vxo���.�.�\��$��V5VM�d7�e���g���B�Oi�G/�'8k��1��?�Ā�E�i�m}66j�"Hs��y��1$���"������,�ǰ'�J:��XD�w�п?G���7�V��i��fj�_V�VG�88�;矷m�w���i���Z�צ���ҧ�Sb4�D�9�Ni�v��Q�P���r�<Uee�,�Aٺ�H���H�V�7�}�!��ϟ��7�4��e���]8\빜�&� yE֩�sJ�|���F��
5[�.������S��?�F�^C��}�����S���� "5�]!�`�(i36���GԸ�����k S���zǣ©���<çI� y?��)(�"����	�	��a��ǣ©��n~�c?Dٿ�O�G������p���r�j�b#!�`�(i3���-���x�fC��T�z���,}l#`�3J�V�h7�mEox�࠿���C��[���ԗ��6%�a¥�����Ј��wfX&|a�#�I7��-5��5Z��N����p$�Q������X;p`�ct�:��RE3z%�u�܆�D:���*=����-��A�sxW�O�,��L��!�`�(i3�nxL�J>tݩ��yI���Ut31�P�V�!�`�(i3&�2�����dv��oTN֢&@��&竷b��"&�N>�`������	�;�ݚ�Н�J�a3mPy��ۊ���<+:0�!�`�(i3�'�al��p�$W�`n\+/��`C!�`�(i3�-���k\�H��bf�?ǉ�=�s�٩�삆-�46_5�(������hy�_�⥳�"_z�Gb��P�!�`�(i3� 䉇o�Mt`�*�S:��IK��<q�\E��0��A��)}��V5VM�d7�e���g���f8���(�:�f,��B�r����n�T���#�-eɤ,��f8���`
 ֢��FE������V��9/RN�]�5'�E�i�m}66j�"Hs��y��1�Y�,��D�.�g3Z�j5�{���������O�A4ZY�j(&
M�K�#7��(ә/��=��K�E��{#6�aAc<�p{סw��"\He�F%�X��k��o������"O��`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��+��%�k<ꬺ��1����t��PЉ�Bk ���E�i�m}66j�"Hs)H��4)�>�|NU�jRV��	��y~��52����� �(㷾���G���Ld�-P�Z:�E����FQ��ݢt\�y~?��
VWk �0D� �B���9���M몴PBoT�G�%LT�:ʽ�fq8*|��@q��=��w��!'|sI��w��,c�A�L'����](p���*<|�����?�������o��C!T*�q���U�h������e�İeR69S�)37J*uV,�������Ŷ;���@��O���Z鎬�������(����c�<Q[j�l���tL��"X��[�����O���q?��0ǽi�*��]�!��	Ǹ�y85��3}�@�7��?E/6 K	����n|#9���t]��\o9%����b3�'���Xw�>�3�J��8�꯮�DES�)37J*uc�A�L'����](p���*R�wX��o�9f1E
�a)�xSsޜ��*ۃ�W�XL�k�T�q�Zl0@���&��c1��v�u�`'s^�`}��AyE0@���&��O��nieu�`'s^�`}��AyE0@���&���� ��
fC��T���i-�̍�{Ф�En7A��^⠻rRV�����K"#o�a�+�wVi:�;��K:SGD@�F��q`E�cvR+v�֐GbH��@hG�������p���Ї�J}�!�`�(i3��`)�pA_g5��pC50����y�;���g���/k�}���X1'1[��o����󖈣���b��famo�C$�{nr���<��W{0`�'vi�K�Ot�td���5
VWk �0'�3=�D�9[8{�n�_ �o��s4k<H��ԇ���M��yr&VxI	�~���A�U� ���_Y�VN�=��Q�>σw�EF�]�`�|��K�z�ix	��GD@�F��q��M��+?�^qk�d	���z�KdL��7�ܥ��2���C�0��(����i����~sv��k�U� ���_'�=�f�J��c:�3d`�|X ����p�IÙ=�H��h�t�����?E/6
� /��4];ˍH�T֟��Bg���j9l��緺4?s�_{X4x�]�V�����TI���0D�Ub��?E/6�ix	��GD@�F��q��M��+?�^qk�d	��e���}����� NM�v#���ޑ؅��FJ��qW8+����PK�k�V�t(]�XnS��z��`��
e�$j�U� ���_V�׍A�M�ſ�lfR	�_�C[��;��6@���sA�U� ���_V�׍A�M�ſ�lfR	�_�C[��;��6`��
e�$j�U� ���_V�׍A�v�֐GbH���x{�:AO����k�*���t�]P؅��FJ��o�C���j��W���Bઢ:g����}� tGD@�F��qW��Ґ�Yj�����T4o64d�k�0*���\�
�=ĭ,Ϸ�@��; G��4?O�!�`�(i3!�`�(i3���D	��U�l>o��|��U�L���� �5�vŞJK��	&Y_��lW��]h�����!�`�(i3"�,�>E����\�v��_�R�G���Fz�Y�b>bb�D���;r�!�`�(i3!�`�(i3�Q�^�y�zL͊�q���?�-���!�`�(i35�K���y��̨!�`�(i3!�`�(i3%Ah�%4
>��XP��ȆS�%�����k����\��>�SS�]�7(��b�!�`�(i3!�`�(i37�ܥ��2���kܪ���*�LNm�k��u��v�Ys�S�)/^;؊���:�6ӰR���&v(𨾤 ���8�TP��k���h�%�F�F=��)E]�� �5�vž�x��&^ɘ �V�	�k�[���!�`�(i3"�,�>E����\�v�T?�7G|`���Fz�����$G���?E/6}�U��!�`�(i3�Q�^�y�zL͊�q��r{= { _m�ڨ�hծ!N�'�y�G