��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�-Q3�Y�K[�J�#.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��9HrbkC �mD�?=j��S
��"C��dKBE7\F���r��C>C�݂�N$��/���	�0���'v6�o~�a�(E
PIU��>v��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&���7�os!w����]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�K�MV}xj\�iW�(� 0�D�A~����p��ؚ�fD�~����pn��-�4ڭ	���
��M!�nz��m��+�q��.���cW)�w�%H�!���Ȗ��h�}�{Sh0�.�	�Z���}fTV����~�hbHp|�P,N��!�Ψ�	�ǳ۱��@�QU3(�R��W�ew2�\�����	x]̍��;����?��|:�-gc�n O�HߵgB�T�V7���p^#����*
��$tU�U>r�O��C��0��ד�̟a�,��I�zb�Z>8��������]�\������������;�kv޶Gl�!��TN0N��\�4�si�W���Y��݅ 0�1���جچB�)oo@���q�&p�`�������N4�$�����(
� �AH�T�t��3��e��ME
^����c�:���0�F@�4%�u�L�r��3�jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��dI�ZS"J��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S)�-E�؟��%H�$��ī�o��<�)�G!�u�����!�M��E��c�W_QL����f�Y!��?��J��(����5�2���[@%����nEA���e�q��'p�@�I�?g�f�P���Z�NCIw4t�iZ]XF�������̅�ԜF���~x�9̺ʆ�In��t����Z����oY��8�b(��,ԯ���gn��s2 �j޽���Ǜ������0Hze���&��J��Vǃ����t���\�W+�[Z��7�ܥ��2����*��>�xn^%��+0�l�R<�jЉ/8y̚[b�0<���E����F��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+"�,�>E���TD���rs�i�jf� l�Ǜ������CyW�f�tR�wX��hs�����n��0�5	x��(�
t��Y�{'%s�:�f~=g(���B��ɓ�~Ҡ	u{ᵿ�����"X��[�d�a�4$�>��68	�-�c�OMe.��xu	�>��l%i�-�}��C˥���6ޭ�@�I��w��,>����C�h�'f RN�By3��<�]�!����M[��Ǣ���ꀍv�ј�"��Z鎬����F�71�B�������%���|g�Y�'���XwI<��f�@O�x�7���9����̠�P\�I������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��9����̠�P\�IL�iײ`��I��'��۟b�/O�=�ͦ����Jg�Z�n��[���M���L�֩T&�eτ�bs��z�h��4h���}둮c_����+�˂߮<u(S2�,̞��>���I�Ūeߦ��R�O�K��ۋ�̞��>���ԜF��O䚥�\�6U����	N�n(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u፦%t6o\N%�4V�H�%'��Ti�ݓ��E�
�oz˸�1�"���q��T�ٮ|�,
���A�;�֋`N��7�j2�ٚC�M�����T�\ ��i3�|)sՀ�|[p2e�F;p�	��2=��h�AԢ�a\��F�dHZ�F�\Ȳ�r�r%)cA�z���a�R�wX��}�
�?���;�/s�1��pғ�vq�\[$Q��
�̞��>���I�Ūe�TU]O�d��g��U-�e,%�0g��Չ3����F�x��&����"���P"G�wk�١��	;q,6KX�#���x.�Knq�z���a�R�wX�ո@����gG��l��`��c%ij��d���0y�	�C�u)�6�3A�)Oq87{�Z�p(���B���ި���������f�T�\ ��i3�|)sՀ�6�S2v:,$��x��f���,(���B��ɓ�~Ҡ	u{ᵿ����2���O��E�%<NR8�b(��D�P�E6�ټ*w2�56kѶ���� �ځ�+W�'/ǎ��+x�q���U��@����gG�K��A��"�,�>E���]�!����w�Հ��pH�:V�^3rdS���n`5�fK���ġC���QK�>;?�ސ�)��1��u�6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>��/���(\w8(�Dt��xjzӝ���I(͂�'�ɳ��!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2�����kv޶Gl7�|g�)��x����E2b�z'hۉ)��d�7�q�hs�����F;p�	��Bf����{_8�Y��=�}�Vݨ��}Dq�f�hzg���5���u�L�x����E2b�z'hۉ)��d�7�q�H�5Bj��@�m�W#�LaX��T.�{_8�Y��=�}�Vݨ��}Dq�f�#��?@�]!�`�(i3��$�\%e!��"� +}0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^�\!�U��0�|�_�mS8<�nVA�ڦ�c4;�E����T��O�T/K���r����KK�+��o��z���	���!^��7���өzW�&��F�u��r��!�`�(i3hzg�����Bf�����;�*�Gx�����}Dq�f��	��x��ݚ�Н����>]&��*j2⎜a�E�Rq���my$�N��o�/���;!�`�(i3���F��O�VA�ڦ�c4KK�+��o��z���	��`�un�&�7���өzW�&��F�u��r��!�`�(i3�⵽2�R�M�Γ�va� ���8#䖭7�j2��S]�_�_��u��r��!�`�(i3��=m緒�!v�/FY��58.��-x�S�ӄz4*�Gx�����}Dq�f�՝� s�#���k$ !�`�(i3�#}�{��7�i'��'DV���b�z'hۉ)��d�7�q�!�`�(i3��Ě�����}Dq�f�HN��R��F F�E̠���y��lD'�ZX^�O�юG�
�0!�`�(i3�⵽2�RH<�2�����3A�)OqO�5���1tSjv�!�`�(i3�#}�{�@�m�W#��58.��-�u:��_xL�[���_>�������Ra])n#���r�����'��o�u:��_x���˃�I��nF���<�W�.�P�	��
�Q�}���%>�rG�@�	����!�`�(i3졾�8 &F;p�	���U�._��ԜF��}�����Hٚ�-����!�`�(i3@�c��F�x��&�"dbnO ��yM�5���%�+� h�ҩ�!�`�(i3��@h G0���˃�I��CH�+�e���;�8w�B!�`�(i3��jVѭ@!�`�(i3H�5Bj��@�m�W#�a�E�Rq���my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp!�`�(i3��z�T�J��	�b��{�Ŧ�4-%$W�Έ�:��Վ�_�!�`�(i3��i�:�3>x�S�ӄz4�XƤ5_�]\1%����_���j�[t�Y81hzg�����U�._�츅��u7rv��$�m��-����!�`�(i3�"�+փIi{�R�$�V��(�iZ`�c!�`�(i3��Ě���ž_�F�$f��_Ub����pT���Ě����>=:9_�a:䩒=]'�Fr��jϤ�Lǀ�v3����t�Xe@�ҹ`����n�3��Z�#}�{��7�i'����Γ��7�i'�N�������`����nU	��b�s�d�1ʮt�u:��_x���˃�I_~h�1g�x�ez8�US�*>�Z����O������6�o8:4��j�V�Z�յ[+8�ϝ�j
������h��`�����y_�mS8<�n�|#HK������ �'����z.��W��t�td���5q�\E��0>�1���sf�e�}s�dKa���z%t��#-ăs��x���ݚ�Н��"� ��.q���f�e�M?��y�!�`�(i3d1E �s�)���Q���3[�u8��a�}�$�&�[.ǣoJ�ҿ�b�K���t��P��l����HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�v�x�w��j�-�]�1�n�cqgF�ht��R����A$�P������5d�	�+�&IiI9�o«IX0F�MТKH�{?��j���A(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R����������A�����q9+t�}�|#HK���؇�M.9�(�����!���|e"�#}�{��9�2�LK7͍��|��W&":����@|����^a�nu4Bޗ��jw�	��!�`�(i3lG%��`��ǚ��ظ
��@�U#�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н��#}�{��9�2�LZ鎬�������(���NTP]�0@�m�W#�	�Ȗ@@��H����NTP]�0�7�i'󻞥O_�Q�؞�(�@~�6Sa쎑�8�h�K7�|g�)���`
�%o�ìzP0�z��:����
�ݚ�Н��]��W�@'����6L״$(�>g�
�:qEp�;�P�t�5����l�� �l�������@+�c_�mS8<�n�ݚ�Н��[�	���"������Aݡٜ�}Dq�f���Ě�����}Dq�f�)�{6�U�����F��O�}�	76�&�� Ӗ�t$�)�vx���Db^3��h�]��w������:?���