��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�4��s�A�|Ԣ��g��B���������'QԵ���
yL��?� �~�ǴW{< &{�!�y�W�BE[��l+ �����)��(�@rD������tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QLi/-�#�~09h�i��I�?g�f�$��P�xZq��t�1�:�Ω��
�/�r}|��ι%9��oGo�Z�J��ݪ��4Z��ʬ�:xK<E<Y@(?udG���q�©����0�w�)�-E������C�x���� �{�7��g��n|��ea�8����U��}�o���#�Pb���ym��+ r���7���?�_�[�htѨݮ�I�?g�f �H�Z��1]���%�Pb���ym��+���uN�YW	��V �T�QT�8���[�htѨݮ�I�?g�f�ja1�n�[�c�/�O��?�;��XC���Y;ҠH�(����5���I�zI.�R7�$��p�S$�&\^�N����{jϾn]��Yk"1/�p�r�w�Sjs����n|��ea�8���B����g��Tݭ�EBÎ6ogN���n|��ea�8����W N��|C��w�Sjs����n|��ea�8��������?9�M�Ч��Dua�\ۂ��Y;ҠH�(����5���ռ�j��I���j{�\^�N����{jϾn]��Yk"1/>���M[�a7Y��0�-\^�N����{jϾn]��Yk"1/��n5R�%�9��o\^�N����{jϾn]��Yk"1/��n5R�%�.��.f\y㔪�_���Y;ҠH�(����5�%���(�-X�Ç�e[�htѨݮ�I�?g�f��m�������d����b���m�+��
J��@��ea�8����U��}�o���#�0��r2�􉢔�S��"���[��ҋI7��-5�B�wj$g�b9���1��]2��2�F�PY~�y�����[�JHn��z���G7���� �����x?����k�c��`��'n�^0op40�zɈ�P�i2s�4<��!I���1��ݥ�U� ���_
`[~&�x/���i� � �	{����0�&�ͭ��|g�Y�'���Xw�f�VHF��>BH<M�z��]���>����CΫa��������-��%Mό���.�DsQ�V�r[%�/��{l�f|�ό���.�q�\E��0�X��?��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A�������Y�r��@IE�U����S8��Ѽm����x?������lC��U�T�\ ��Tǯ�!���#;r�����S��I�?g�f�,�� zr����$l2�W�K��q��"�$"�N�p��G_�(����5���&<˴m���q~�i��Z�NCIw4t�iZ]XF�������̻9Cd��醚/	�IJHn��z���z�O҈�]V�H7'�R�^Ƒ�� ���3�ҺIÙ=�H<z,Ҽ&�z~~�Y_" �g8YwU��֜��3JHn��z�Sp�}�f��]7K�6����it	�T�=��?JHn��z�ڒ�/;^�/���i� � �	{����0�&�ͭ�E����F��j��\w��0]Y��
�iC�E����F��j��\w��0]�\�LtF��E����F��j��\w��0]EOJ�uxm�3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��D�@�Y�4��j�O$� �P�%.^F�	��lC��U�T�\ ���A�����
����Ř]2�y�Z鎬�������(������t�\~ �g8Yw�5�%]���a(􆿳�ؖ��d�I�� �:&�� VU+I��vMb��s��Yk"1/]���!E�TU"��JH3#��Aq��:9�+�m��+ r���7�����|]�Xy8��;6aJVlO/8֩]=$���4�+|'�kP�?qNzL͊�q��UG�s���w¹��<d���<
DN��b9���j}8o{:�d�}Bȱ��U�p�[��i��i�����8�TPF�� g���t�&_���9��E����F�'n�^0o��ҕƦn+0�l�R<�q��f�}��?��[�<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����(��eظ��7�
BcyMu򔲊'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5��6��	���`y����ꢤ�Og�?�#B,�Ң�{l�f|�m�jp=�>��o�
�v�ξ����LUG���>��Oޏ��F˯�+)�"j���b7|#9���{k�h�++k&v�Iz7G#+�ǚ'b�t	�U���C��O]r�<Uee�,��3�L���&Ã�M�R�^Ƒ�Өg��U-�eaԗ5��C�W�T ��x���� �+��T�����h�6ؖ� onc b�Vg�x���� �+��T�����h�6ؖ�{��^�
r��4�3dY�-�nC/$jQ߰�H�M��RV!�`�(i3U��֜��3����C��n����e;��}Dq�f�S^�1���yد�9����)h����M��%�p@��\ NhJ���/�UI��?X�c"`.� �#�i0�[X�b\gA�[3�.!�`�(i3�=��?Q���n�;�X_y�F�!�`�(i3�{d��L����Oq0}�+�]}wӭ����?�+,���iVA�ڦ�c4���^���.�c��><�$�z�)
ԏ�.T٢ߡ[�1�g�=��2U�u�H
(����7S��Ro8�ih���
�e�~w�!�`�(i3!�`�(i3!�`�(i3!�`�(i35K�,<J��.� �#�i�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3ԁ�42����t|��z�W87"�o��ѾJJ�����	.l�@{���e����P];�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�-��\���7ȡ�/�!ҔkmB����I��%�)��!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�����-VL(;�D��g�FBZbQH8�I�we3��r^�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3m�z��P���ڞ��3*�f՗h�Vdoq�M辙�
so��j�!�`�(i3!�`�(i3!�`�(i3!�`�(i3MX����C���7}�jA�� <LS�ʌ���p5B���� �o�X�S��Ǵ��BE���Kt�I�ZMz��v�N`Z�NYUO��z�W87"�o�j'��y�?&�2�����B�X
d�E U�V|���hy�|�ր9�j���B���7�F����|��p+E��%>zcbp��'��}Dq�f�4��d�X��H���z{<���낌״$(�>g�!�`�(i3)�{6�U����/��w�=�J�5x������l����4�n���xǊ��T�3,R�^Ƒ�ӳt&:���aCPW�����8fDs;ly��\%�0�9&،{"�Lެ�k<�Lơ��*T�Z|{�0z�cULD�vO��|��!��5:A�8���/�l|�*"k���(ӈ���m�r�������Ȋ�?�Qs5��uYl���#Kv���:1�#���FT����fK6�L+�.8%�����dN�<@Iv��nt=:�rl��7�L�{	�����Wm�0b��"B��$%eqq�\L$�����//��kOTm�ڨ�hծ<�6�Q=a��	�sǡ �w�;>cbp��'@
9��yž
�I�>y�t&:���aCPW�����8fDs;ly��\%���y��lDJ�z`_�z^9;����l����4�e�kzP��}Dq�f�)�{6�U������ł�me":l�n(��̓iq�����f-���bX+D���0�7a
��r��X~L��U���N���{_8�Y��n3��v2!�`�(i3�ǽbI�͎DX��,�6�HaDl��+BY��9�)(����������qϛ�M~!�`�(i3�ˇ�h��]�Hlu�����}Dq�f�4ﲐ�if���ٷ����
t��{<���낌)P<�ܓ�Y��'T���+\��.��4��!%���Kv���ft�s� uƍ2���l�A�����2>�>���v�|��z'���Xw�����C��ݚ�Н����v�gY�����Iꑤߎ��J���T���b+}y[���S�fh�����0�T<9 =��9�j���B]��>��y�(�Tl��z^9/�~��	��D܂�A�N�p��G_�(����5��x���|�:S�Q�[����g�� b�Vg�x���� �+��T��/o��إ�8p	�rh5���Z=%��0��r2�􉢔�S����j�}�I/��=��K��䘾is�%Ah�%4
>��XP���G\p���q��Q��O�بeD�I��[7�d|���XP���5�%cOL��5��Dz��!�`�(i3%Ah�%4
>��XP���4֔ʽ�I7��-5�B�wj$g%Ah�%4
>��XP��Ȩ�wl��h�Vx�%L��]n�� ���3�ҺIÙ=�H<z,Ҽ&W����vcy��<
DN��Q�^�y�zL͊�q��ø�B3^�MNM(�n��1�Z���=�i��i���'n�^0og��jU�U��2��̪
)\Y��"�,�>E��4];ˍH�F�n�ܱ�7̧�����A�����y������i��E����F���8�TP��������ERF�G{؍��R��j�.(Wx*��|��pe���b������5	���]���>����C�h�'f R!�`�(i3��|g�Y�'���Xw�E�i�m}6�B�r���E����F��j��\w��0]EOJ�uxm�3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��ct�:��RE��W��_�ړ8���/��^����r��H�+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�H�NI�:7�N�5�%]���a(􆿳����^��+��%�k<�6��w������
L'���Xw s4S�'�i��`�z6/������,���eFz����zf�U����z~��6��	�\�HP@�a%=dϖ�i��F����U��:9�+�m��+��jTʱ�8F0_H��w�Sjs���h���G!��:9�+�m��+��jTʱ�:W���	�)�0�lOw�Sjs���1}Kط��4q�������o)�]r k�|6�8�����JHn��z�Sp�}�f8֩]=$���� ����H�ʱˡ �ϭRoF�'n�^0o�pJ1����^�F��M֋)�[���6�E����F�'n�^0o<H�-��*����Kp&�@���k���E����F�'n�^0op40�zɈ,[�=·j�U��֜��3"�,�>E����\�vņ�Q�]����O���R�^Ƒ��!�`�(i3JHn��z�æ<C}�E�먾�� �Y�7#�xI��]n���b9���e�ʼe Ej޽����3i�z6���������D	��U�l>o��|���/Y$�cA�\.�
��ڃ�"�!�`�(i37�ܥ��2��
[���p�� +@����wF4��0[����	��N�Ae�#����ꀍ!�`�(i3c��Et��q���U����?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-�|�)՜�4!�`�(i3v�ј�"��Z鎬����(��eظ�_--���g&e�l�����-��%Mm�jp=�>��o�
�v�ξ������ei]��fM?R�^Ƒ����"X��[��Q[R�7W����GS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l����G<�e��
T�v��1���6��	���`y�����o<|O��%�ꤸ���|K��h��?�w-�%��p�i7GeY�+��%�k<�6��w������
L'���Xw�j�7���i�_:���5�%]���a(􆿳�te�"���$+�uB;y�L�6yd(��(�
t��Y�{'%s�[�&B�踫g(�r�2�������l혡�[�����ݪ���CyW�f�t<|����faՊJ�	��D܂�A�N�p��G_�(����5���I�zI.�R7�$��p�S$�&�u���k�ȻD�ou�*Y x�S��q�©��ല���?�;��XC�,�-fce��,\ަ�It�k\,آ(&l������ nU�IÙ=�HF���m¡p~z�r,i��i���'n�^0o<H�-��*����Kp&�@���k��JHn��z�_c)���8�+�p}>&�&i�A ��E+���XP��Ȩ�wl��h�d�uY�ة�ʐx�?�'n�^0o4M,������2��̪
)\Y��7�ܥ��2��
[���p? E%n�/���i� � �	{����0�&�ͭ!�`�(i3N�By3��<�]�!����M[��Ǣk/�z�xEQ!�`�(i3c��Et��q���U�&��GE<�!�`�(i3Y%T��BPe.��xu	�>��l%i�-��TBd��pS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l������\�*P�I7��-5��6��	���`y���db�\EX@�/�M^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'"�C�ף�;�¬pX��g��U-�e�,���6+�+�uB;y�L�6yd(��(�
t��Y�{'%s�[�&B�踫g(�r� k�|6�8j��RO�I�1�Z���=�"j���b7xY�J��ev�mS��0�
���)�*Y x�S��q�©��ല���?�;��XC��z���ْ5
�8��1�:�Ω� C�`N��D���ÿ0�^��pZ�NCIw4t�iZ]XF�������̘�иܖ��i (LW4�'n�^0o_
-��[�b�ӝ5�T�@���k��jݭ�F���L�D��6S^*?�z�̒h��l0��F��j�mV��5fj޽���Ǜ������(���{�OF8<z,Ҽ&��v��z�N��������\�v�C��=x��ҷ��.G�U�����\�� jZ^��ecT^�`T�W�88�;矷±�sR�{F3�_� ��"����5'C��[����N�pS��Y���8�TP��Vch˪��/h�h��=���Q�n���{�)w�<�_N��}��|��hLbLrB(��\G�Y����-�,�.y���,�x��#��]����������ݹ�0�����иܖ��+V.���A�sxW�O���lC��U�T�\ ���A����jsrCm�k/
�ȡ>I��w��,�������ݹ�0�����иܖ��+V.���w¹��<d���lC��U�T�\ ��+�_0c �ۧ2���{�ҋX����>��l%i�-̇i�d�?���{l�f|�ό���.ӳ�
�	?�<7Ê7�E�4'���XwI<��f���nܰ��ْ5
�8��1�:�Ω� C�`N��D���ÿ0�^��p b�Vg�x���� �+��T��/o��إP�e`b�T=am�����/�����,��B	hI�ˋ���p�ϵ�DE�U���w5#��1���XP�����<��F�r�f�t?�1J&�|D�e�!��L�D��6S�]V�H7'�R�^Ƒ�ӥ�e%)>�Z��&��J��Vǃ���O�4ۤ�`�	��B�f�\�kA�/����<.+6J!�t���\�Ws��l=�L؅��FJ��G��k���؍��R��j�.(Wx*9��?xs���}�ڍ䢝{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�ս��Mڷ����}�ڍ䢝{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�Ռꢤ�Og�?�e����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+�+�uB;y����f�O�]�!��M8���	D%*`�u��,�Aٺ�Ha(􆿳�56�P��/�5�%]���a(􆿳�ټ*w2�56a��p��)��{l�f|�ό���.�4%6� �77Ê7�E�4'���Xw�f�VHF��>BH<M�z�]�!����M[��Ǣ�:��6�J�ҋX����>��l%i�-�|�)՜�4��{l�f|�(0̈��N�faՊJ�	��D܂�A�N�p��G_�(����5���.�^�9��ǘ^�?�;��XC��z���ْ5
�8��1�:�Ω�>���U�_�4�0S�����x�/�����,��B	hI�ˋ��b�ӝ5�T����-N�ʆ�In��t��GAџV��2��̪U��֜��3jݭ�F����QI�D/����ʊv.s/�B{�o
�_ q1j�iϳ��溂�U~܎VV��EfVNNwK35������8�TP��Vcht$W�<	)��j)yc�n�.�_�t�7�ܥ��2�΂��F�V��Q�S���>³��w�[��C��=]A��O�T=�4e=��-������yM�&B��S��+0�l�R<�q��f�}���D)���o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y������q��w�J;QPטeS�)37J*uc�A�L'R�o�����5�%]���a(􆿳�ټ*w2�56�[b�0<����|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<� ��i)Y�I��w��,c�A�L'��!�a��5�%]���a(􆿳�ټ*w2�56�Aɀ��{l�f|�ό���.��_F�k-�7Ê7�E�4'���Xw�E�i�m}6*�3���f�]�!���D��L#�jAY4 mv���S��I�?g�f��Qө}�8o�C���7I�����u���k�ȻD�ou�*Y x�S��q�©�����<��������/�����,��B	hI�ˋ��b�ӝ5�T�@���k�փ��㛋��X���`��.�̀�I7��-5?�1J&�|D�e�!���QI�D/����ʊv.s/�B{�o
�Y-�E�f�}�=Ll�����,۽���}i�@�5�}�]���x�]�V��7��_��T��!e����\G�Y�)��Y櫧�7*9uu"�,�>E��<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9���[�t��#���j;9ekN�By3��<Z鎬�������(���P����ˮ��lC��U�T�\ ��+�_0c �Q�P��
S��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+�����
L'���Xw�j�7��ct�:��RE��W��_�ړ8���/�z&v��\��t������S�)37J*u>����C�/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�ЂDa��(O�J,���Z鎬����F�71�B��O1��m<S�)37J*u�񁫴}2;9�".<�x���� �+��T����oGo�Z�������--�p�,X|g5�GX�����S��I�?g�f��Qө}�_g�?�H���w�1K�E�\��Y�ea�;y� ����t��A�sxW�O�k�c��`��Z�>)��`�U+�PA����Kp&����-N�ʆ�In��t��Q�]���h�S{�5��lW0�±�sR�{F3�_� ��"����5'C��[����Q�n���{�)w�<�_N���i��I<��fҾ��9�ǈ�5�G
m��u��N��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�D�+���8�<��z��}�0z�cUL�n����4���á�~O�"j���b7���Øfq�\E��0�ŭ�����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��Pc�Xe��TD���rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0���-n�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�eן�-�Q�Z/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�ЂDa��(O�J,���Z鎬����F�71�B��O1��m<S�)37J*u�񁫴}2;9�".<�x���� �+��T����oGo�Z�K����ހ d���j�޺�5%��m�+��
J��@��ea�8�����B}rs4��������b�1}Kط��4q�����Pq�=6����+� ±�sR�{F3�_� ��"����5'��иܖ��i (LW4�'n�^0o�pJ1���ٵ���Kp&����-N���\�vņ�Q�]�ޔiyV�[R�^Ƒ���b9���j}8o{:��͹ ��1�Z���=�A ��E+���XP������,��=�$�ЭU����z~��;ε��IÙ=�HF���m¡f�Nd+l�Yҽ֗��[7�d|���XP���|t�N�9������e����y
 <JHn��z���G7������=�A���ۖ��S�<Ԣ�JHn��z���o�K�Dd�KPZ���<om���[7�d|���XP���nN#⦵���Օ��qvdЧ^{�j�b9����4�6�t�8֩]=$�����k!�\Z��K���b9����4�6�t�8֩]=$�����k!��V�_g�JHn��z���G7�����(��q�
�Bk�i�����B�[7�d|���XP����G�u��ߡH�� �Y�Fck
���/d�s��p��'n�^0o���˟y�A�o��d����O�]�A( ����_ֲ��mŹ�[�g�DPp�A�h��+FeA'�u���.���hGD@�F��q&�G"�2���k4�͹ ��qC��~�;ϔW���1��ݥ�U� ���_�g)�X�:�G�
f�V�5t��\�H��/Sg޶��g�R6ӸJHn��z�1��-�\{]��ˀ.�� ��H}ة2�IÙ=�H��'�PD�C��[���ԍ�7�"�����=���aw��Y�ڪ,[�=·j�C��[���ԍ�7�"�����=���aw��Y�ڪ���E_����+�+#B��1��ݥ�U� ���_?�(����۫wH�HͶ�t����oD�c=p�1n2�I�U� ���_-�"p�)KCs 3�:�}��oFkZ�U� ���_������yM�&B��S��+0�l�R<�q��f�}��Gظ0����Y%T��BPe.��xu	�>��l%i�-�M�g�����E����F��j��\w��0]%��C���M��cg�P��-��%Mό���.�y@�,�Y\��_'�pfn� N�RZ鎬�������(���{� c*v�T����1ܚhU_��_��Cҷ��e�ˇ�h��<�W�.�P�	��
�Q�}�˩��*���"B��$I��w��,>����CηxmQ,ۘS�����E��@IE�U��>��l%i�-�[b�0<���E����F��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���EOJ�uxm�H/t��)��-��%M�:2QYeƈ)P<�ܓ�Y{k�h�+"�,�>E���TD���rs�i��~Ȃ�D�1�Z���=�"j���b7|#9���|�au�(Z��I�V�~��TD���rs�i����ej1W��Mw���1�Z���=�"j���b7xY�J��ev�mS��0�
���)�*Y x�S��q�©��7��#!l'���h�W�ӝ:X�{!�'R�{ɟ=:�ْ5
�8��1�:�Ω�[@�qR�� ����L�Y�͋�<Ct�z&��ÃlO ܅d:`q裸�Pe�E"��B�wj$g>���'hZ���溂�U~܎VV����M����3��~ !�`�(i3JHn��z�����͉�]V�H7'�R�^Ƒ��!�`�(i3%Ah�%4
>��XP��Ȩ�wl��h�Vx�%L��]n��"�,�>E����\�vņ�Q�]�ޝ��(��U��֜��3!�`�(i3%Ah�%4
>��XP������,��=�$�ЭU����z~��3�Q��\�v�T?�7G|`�LEƒ�$�f���-A�¤�x.�Knq��u*K6H0�T��:GҚJ<�(J�.ᬵy���gP!%�d�Q�^�y�zL͊�q��1�KB|1<\��M���R��ӟ-�������i�JHn��z���G7�����o)�]rx�y�Zgl�q	���%Ah�%4
>��XP�����Յ�(�����O��86�E����F�'n�^0o���˟yD:�����,��R�c������i��a�\����H�:"�\��}i�@�5�}�]���!�`�(i3���+�J��U<o^.K�}��HwL�X�+�p}f�~�ڳk+�[Z�����+�J��U<o^.K�}��HwL�XArߟьvb^:�x���1)fd�vĻ���+�J��U<o^.K�}� c�2��`?iRPsf�Nd+l�Yҽ֗��[7�d|���XP���&��@2�G��&1���Q�~G%2����D	��U�l>o��|��v���?�5�h�I�nI�`���1�Z������\ ���+�J��U<o^.K�}26U� �K%U���?��>7�M�Fri�u�q��k�ʆ-�H\���IÙ=�H��'�PD�,Y�o�a�gf{}#k��Ȟ�����i�U�4��X�Ặ��Ϊ�Q� ~�����(��q�
�Bk�i�����B�[7�d|���XP����G�u��ߡH�� �Y�Fck
���/d�s��p��'n�^0o���˟y{,�
w��|ݔ�3�5�}�]���7�ܥ��2��Э�)P�q���Ì �&�k��>���c��d�|ݔ�3�5�}�]���7�ܥ��2��Э�)P�q���Ìݣؤ	����2��̪
)\Y��!�`�(i3���D	��U�l>o��|���/Y$�cA�\.�
��ڃ�"�!�`�(i3���+�J��U<o^.K�}�������ɰ�͝�e>����C8����̇i�d�?��E����F��j��\w��0]Y��
�iC"�,�>E����-��%Mό���.��6[��u�V�<�nbBIc��Et��q���U��^L��6�}�%b�CGފ����]�!��	Ǹ�y85����!��K|�d�MHOm�<G2s�%�8���/�l|�*"k���(ӈ���m�r����h��eZ�����E��@IE�U��>��l%i�-i��H�p�E����F7G#+��\w��0][�л���7"�,�>E����-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0</���/�u��(�
t��Y�{'%s:3���5C�ݪ���CyW�f�tR�wX��hs�����n��0�5	x��(�
t��Y�{'%s�h�v���&���$S�ݪ���CyW�f�t<|����faՊJ�	��D܂�A�N�p��G_�(����5�%���(�-X�Ç�e8����Bp� VU+I��vMb��s��Yk"1/+���鷦:`�'ࢯ�,�-fce��,\ަ�ItK�1�֎TW������������i�l0��F��jT�����N��3w:��ݪ�򈟞�����i�%Ah�%4
>��XP������,��=�$�ЭU����z~��;ε��IÙ=�H:t@���8����̇i�d�?��E����F��j��\w��0]Y��
�iC"�,�>E����-��%Mό���.��6[��u�V�<�nbBIc��Et��q���U��X�=)�H�7M��񇬦���
L'���Xw��+x�r�2�6�d�f�]2�y�Z鎬����(��eظ�=�tneX N�By3��<�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+�� }'�8�������5	���]����,�JL���ƍ2���l�\.�l����"B��$I��w��,c�A�L'z��0N�7;�¬pX��g��U-�e�,���6+��kv޶Glbq�Z��T�I��w��,c�A�L'�b��9X�T��&��;�¬pX��g��U-�eaԗ5��C�Q�$�k\_x���� �+��T���O'�lR�����|7�:X�{!�'Z6:�q�_�x���� �+��T���O'�lR�ܓ>��iכ���������N]�Xy8��;6aJVlO/8֩]=$���GZ>.�0�[7�d|���XP���<����k�|ct�:��RE��Ok��@zL͊�q���Vǃ�����������-N���\�vņ�Q�]�ޝ��(��U��֜��3�b9���с�'sIP���1>y���Mw���1�Z���=���u*K6HT�����N��|�P~)x�?{���x.�Knq��u*K6H�q	k���AGҚJ<�(J�.ᬵy���,kM:�yzL͊�q���bF�����M���R��ӟ-��[7�d|���XP���|t�N�9���r�&U������G|M��[7�d|���XP����A�\�n���~�����G�٘�Q�q �&���M���HaU$kX��� nU�IÙ=�HF���m¡A�h��+Fen����9��#�B�sYC��\�v��_�R�G�$����{v��G�K$xE�p4rqG7��u*K6H �i7�sp>��%��H��5[�����q�_�N�6�Ặ��Ϊ�Q� ~�����(��q�
�Bk�i�E?�xu����ma��u��ۯi\�q���Ì �&�k��>���c��d�|ݔ�3�5�}�]���x�]�V�����Ү��`�+S�p��ͷQ�X��9Wp��� ���U��7�ܥ��2�\Z�ؿH�jGjh�rO-�<i���A���U��7�ܥ��2� �2 ��գM��b���=|-�e1|E�A�2����ma��7I�����;�h�]�6�F)=�5�e$�m�w�3�a8&N C^�A�����y��7�"�����=���a,+$\�M���j��"n+0�l�R<�q��f�}��Gظ0����Y%T��BPe.��xu	�>��l%i�-�M�g�����E����F��j��\w��0]%��C���M��cg�P��-��%Mό���.�y@�,�Y\��_'�pfn� N�RZ鎬�������(���{� c*v�T����1ܚhU_��_��Cҷ��e�ˇ�h��<�W�.�P�	��
�Q�}�˩��*���"B��$I��w��,>����CηxmQ,ۘS�����E��@IE�U��>��l%i�-�[b�0<���E����F��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9�����E?��� �	p�	��|g�Y�'���Xw�����C����H��?�0q5;�F�{k�h�+"�,�>E���TD���rs�i��~Ȃ�D�1�Z���=�"j���b7|#9���|�au�(Z��I�V�~��TD���rs�i����ej1W��Mw���1�Z���=�"j���b7xY�J��ev�mS��0�
���)�*Y x�S��q�©��7��#!l'����z��d��o�vC��h�:EO����S6]Z��K`��$�dea�8���A��>s>;�u���k!N�'�y�G