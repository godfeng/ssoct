��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����Q%b<Y�D �c�=0N���6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,�Q��Կj��_�L��o¸���Pq����w�Y��k��ı����~K�%��w�Sjs���N<��;��� B]�pE���	x]̃Dj#^Da����M�ٲ��9ߪ�
�M��ļz����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��� ��|4�)�����|�1R�_ߥ�]��4�:j�l�,9���U�/�kl�F�..����+U�	��  �ݘ��`��О������/��^���4!����Y�f��a�Z��Vv�c
����7(�(���2���oK���j��J"/��B������0�M�be8Wg��5F��(	��������E2ܠ�􋒥)��Hi+�3��������*��pcg'���>;#�|����W���~=�L��/f�G P=PLF�Q$�Cte~t�:>��Fr��x�|Y4Z�S��N����PT]e�5{����k`�o�I\\+�����p���Rd!rf�AO]|�]zz���l��׎o�| �mHbw3v7�9��t�,�;��Z,z�eq.��B�0�����'m�b_�V\Xո}3�^<�^&2��m�/�S3 <;�:�d���j14�"ų��K��f��������[|Y��?{�Ac��2<Fl�Ř#1[�3� �������Q��[�x��K�h90�j�����JN�`E�p���QJ��m�ק��-��X����?�ĻY
���+}��������W`&c�'N�j�Y����<\by�5��4��g�:��U��ob)^bK���Ťr��urM08�����x6<9�P�طPӢۼv�^a*j�x������MK9(?��l�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
2,w���~�?|�[_wȵ�e�kY��Y+]��=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+���c�W_QL�ѬL�1m��+Y#_WӢۉ���2=�l�������+rb��'f�ٵ�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/ri�y�!�3]o��in�m��+�<4��ˌ�ň��h��֑�/6K�RZ�NCIw4�ea�;y� h[M	:$U��֜��3!�`�(i3�a�\����9�	��%�	��El5]4 :��	�φ�F��F\��\�vňu�,�s���ǁ��f6�=��? ���3�ҺIÙ=�H|�&��@k�C�H�Lg��DW�3Y��P4�4GJS�x�9�f��!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDp��<d>ARp�W��9g�Z��b,���Q���x�#r���F7����A��=O���[7�d|���XP���fB	�aR�vbR�K��������A( ����_ֲ��mŹ�[�g�DPp��־5�9\��]���#�ڊ<?@Pʶ=�����|#P����τq"�;�.ʧ)ߞ{�l?�I�� 2�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���W��Ȑ:4wh GqH�tU���L��a�h&gR� �ұ!�`�(i37�ܥ��2��
[���p�� +@���x�j6:mU9����u������i�7�ܥ��2����*��5�V��On+0�l�R<�Q�(*w��k/�z�xEQ!�`�(i3c��Et��q���U�ЂDa��(���o�d�Y%T��BPe.��xu	�>��l%i�-Kp(����2�����VcƮ��.J� ���rqϟ<�^�5��q�\E��0!�`�(i3�"B��$I��w��,c�A�L'�����CyW�f�tR�wX���D������Ҷ����S"�f'�gܜ�]����$u$Yo�K�f�NF��D�,�H���D�Ͱ�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3+0$�oI�K&������f��Gm/s
9��
!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� �JB��7C%��ـ��Ϝ���}b�z|w:R��D������^́|�A�"B��$I��w��,�$u$Yo�K����$h������7ÎƖ�"k@:G�!D2W��!�`�(i3!�`�(i3!�`�(i3!�`�(i3M�8Z�XPt(o���xn�q�+��B	cB��!3C�4M/�S��ݡ��1��Yl���#�]�!��	Ǹ�y85�����F�>Г�����g�>x���φ��0�jS�X(5��+��1Ld��&KG!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�O� ��G�P�U��Q�@N�
ǹ� �Z8��
��k�\�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�������F�
ob�@<:�Z1/�ve���� �O�DC2+E����[�`S��|���Yl���#�]�!��3{ح���D��r'ىnX�n>���{�$�˽�L��"k@:G�pP_��G*!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л���O)T�;e���p�����"��3v�}&���s+"�t��gu<�����E��@IE�U��`�-9v��"�����B���>��d�b!��u�4�����7J|et����$!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD���bxA�����|*>i�ܻ��`��_���¯��M��.D�+���42�����Vc��;�?�F%I�����9k!����N�1�Ð
�����=�	�/�2���TD��-�`��8�45�V��-����D��ܒp�@OM.Ir��������ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��7��"zF�e{iʖ.gX���4�d�W�� ��lp������e�D.7�5���S)���-��%Mό���.�^	QW�Q!r�!���;�����5	���]���c�A�L'�����CyW�f�tR�wX��^	QW�Q!r�q� P������5	���]����,�JL���ƍ2���l��K��I/� �����c��Et�p�VU��Jm�QA�Q* ^	QW�Q!r~$�}>���*E9��?��]���c�A�L' ��a���1;Z�减o�ygJ�ƃ/���R�y�� �d!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD��kط����;d�)���l4`��뽣e΋���B�Ӑ%=dϖ�i�@O�x�7�k�ZV"���:��#tC������s��Z����g����<ë��r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+�<4��ˌ�ň��h��֑�/6K�RZ�NCIw4��g�,P�n�U���q�
@�<[n^/���$�G[��&�v��%eP�� ����Og�r�B��9i��TCl�`4_r�Hl��T�e��r��O5k�I�KO��&�o��E�
�(�����;v�BI�ڵ�  $E�ʘ��`�78>�S�=":9�˭;{o���z�r&sq�dט�w�� �RNKr�ɢ�"u�����Y���4�'n�^0o�'vX[��vW4��`���\(ܪ����)M��dט�w��׺8|MW���0o�_o��E����F���8�TP�M��=�&&ĕ^$&��Z|�W3���U���֍z����I��'�^�~����U 1�|1#��Z�����XP�����C��`�'��q�cY��O���vIH2l}�{rcKE#��_/�}_�7��
�+�0]��$�'�k�H��Ѝ���eئ�=ߙ�@�1�˓JHn��z���|��Aו{$�3~��E/2L#�A%��@���_����'m�|g�~p!ۓ��������-���$��Xo��� ���Lk�=�א=ͼ�\�v��� ��o�g�&�0m��Dػ@3�q��f�#��@�RO	�]�ْ�E���$���ş�'�F'�#aZ��qA�E�������D��ɍ��/f�6's���ZBi�mR!.<ή�$	�:-!@xNr��졾�gD��ɍ�ٷ^��o�9p�̺���}�
�?��hҜ����_ɵ@���Q]� _ό���.��7�b����U�m#j[�ߏ�����e��Ek�Z鎬�������*�n�B��DP֞ ��o�;Ĕ4(�U�w�7s�9���o>��l%i�-�����bp�}���1�#��d_7s�9���o>��l%i�-ݓ��E�d�>��W����}���7s�9���o>��l%i�-ݓ��E�F��6�!�`�(i3q��T��|����5��"u�����2����/�g��U-�e,%�0g���j���'l/7w|] ���}N�#�ڊ<?@���,D�d^�-Z���D�kJ���i�#Ѻ'���Xw���,Dߔ��� �3y���(���G
'���Xwd�n]N�/��A����Q[R�7}ϼ 8����Ƀ�?PA�ʻ�(%�7s�9���o��S8�P?_������`y����˞�Bx$�Z�0�]Z����"�,�>E���]�!����w�Հ�>Vۉ�!=5.B������1�U���]�!����w�Հ�>Vۉ�!���ևA��1�U���]�!���e��Ƥ5�e`��94\%��t�E�`JcU�n`5�fK�\w��0]7��"=���Li�ҠG�����зq8�Ј'���Xw%������d](ùy�;�b9����U_�+Xٕ?�0V4 :��	���+!_\�/�@����gG7�6>ᙇ��5ǗcV�j���+�J���q���U��@����gGT��+𦊢��^�v����+�J���q���U��@����gGT��+𦊢BwH4��~��E����FZ鎬�������*�n�B�E �����VF�˷������N}�d�٣���N N�S��E ���� ��M�#!�`�(i3�d�٣���o��D���/h�5�G�G�B�+2����_͍��n`5�fK�\w��0]7��"=���.ZQ�*�3���g����+�J���q���U��@����gG�8��y�lت�S^J�Z�d�٣���N N�S�D[��+s�ceb�)ZF�1����U'�q���U��x�6�u�Xf��@;��,i ���}�CU�+vό���.� ��h���0�`x�֒���\��n`5�fK�\w��0]}�
�?�^���+| �g'#0fO'���Xw���,D���6}�"���@$��]�!��!�r�C|T�He�-�cW8�8J�|9���7Z��7s�9���o>��l%i�-He�-�c��3E M0���oww�7s�9���o>��l%i�-He�-�c��d��]�QS���c,�]�!��	Ǹ�y85�B���0���u����g�&�0m�7���r���ˇ��$�'	�|#9���7��"=��|�w��DK����$������+�J���q���U��˞�Bx�T:���V��pu7����E����FZ鎬�������(���Jם����"X��[��Q[R�7��B�D�F ݰM�_�G]�;o�� ��7s�9���o��S8��y�)xʔ���6��	���`y����@����gG2^o�!���!�qg_�S�
ut�q���U��@����gG2^o�!���!�qgޡ.pz�Lۘq���U��@����gG�5�3�������kO���+�J���q���U��@����gG�5�3������� +���+�J���q���U��@����gG��d5C[�[40����x���+�J��Y�{'%s�Ǹ2���$�mo�6L�g��U-�e,%�0g��ա�a�e56<#λ��$S���c,�]�!��	Ǹ�y85��3}�@�7~WGS��yB|#9���b!��u����ꀍ!�`�(i3�n`5�fK���ġC���}�
�?�U�07�:��=����h��Q��ۆ٘�� ��`t�A~�@����gG������PȮ۔��5�'v�]��������,L�k��V�4�I����"���XmIOñQ��]��]�!����w�Հ�ꓱ�ҥ ���_�,)ȍHK�O��ӣ��q���U��˞�Bx�)׺����xV�(0�8����C�q���U��@����gG�uWb�'8�B�>�zViWS���
^-#"�㼱ΛwV^(�=#v�PriDJU�kTv>�*���i��k�ȓ�iӚ/����C=+f��!�qg�-��h��Uo�A������u\\�~�<��W��j�[O����k$ !�`�(i3!�`�(i3��qTvwN1��\���S)G�6�!~���x�����뒋N, �c����w�����\���S)"�x�H��H�2^�/3!�`�(i3!�`�(i3?Q�@X>#��ŕpO"
P���@}�QlS��3�LIhgN�,�	ܷ�4D�P�>�s�,�H;��|B
y�3~;�>�Fr���A�qIp��K�+}
��.ό���.�d=��¾ȼ^	QW�Q!r~$�}>���/�k�2�������Px"S�#�dń��,�HK�Ƀ�?PA�g�+C��s�ܮ2�k���xw�F��~��;��x[�2�х2�w���㔍�p�׃tUo�A���K��I/N#~8"�Z�q�A��Д	���QC��{
B)U@ڸR9�)L*k������k$ !�`�(i3!�`�(i3���%��Y�Z����r����%6��ڥ����Ⱦ^�����4�M/*�3�2��
 JSV`t�j�O��[��o}��~�f�����k$ !�`�(i3?Q�@X>#�J֎GJ�.��K����-��h�r���t�T��4c�� n�ƫ�}<�[��l�,�m��?]M�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3s� ��<C
�M����G�k�a�`^�Ad0�|��'N[��l�,#̋�X��Ad�G}%����3f�B7�Q�+ż٧��>Y��߆NU�
{�~j9}^p�t|�7Ԝ7(u�!�`�(i3@��]V8ml�i��- �!�`�(i3�B�+2��;�P����|e"�H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3����3��[<�m��I�՝� s�#���k$ ����l��T���ӄ��!�qg[���**���k� �ԬQ���Kͽ<\��1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=I�^$D���������P�íN=]a��o���H�RtV�^!�`�(i3�<@���ل=����h���}�%Dܭ��}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/���%s����K!�`�(i3�̢k���������P�꠼*d�m�d��-��!duP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���QCH�9#G�>������
�:qEp'{w#/ B!�`�(i3h5���=�t���_j����ۈnp� p��@���!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �(*�O�q?qV�s�� �ݚ�Н�
̛�]���n���G΂��b+}y[!�`�(i3]���\�x8���D�kJe���N�ScM?��y�!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3��jVѭ@!�`�(i3,�˳�*C[��l�,t���H[W?��	P �a��e�D.7�q���f�e�&�U��f�!�`�(i3����&��r��졾�g�Y������y�!�`�(i3�߆�p�h�T���ӄ��!�qg[���**���k� �ԬQ����5��t�1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=b~*��s�������P�íN=]8k��.ͥ�H�RtV�^!�`�(i3�<@���ل=����h�]
���7Ϝ�}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��OEʨ�`N/������&G!�`�(i3�7����������EN.74/�������yr�!�`�(i3�����!�`�(i3�7����������EN.74/���g!�%=F�=!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	������6���WW	�Ec�&U�)j�S���vo� ��M�#'�^�����ݚ�Н����g!h!����e_�g�+C��sG��Hb� h�ҩι�+�t2��Lq��QF[��f�\%�,�F��P��}Dq�f��	��x��ݚ�Н��H�����K��I/z�
1���;��J����
%�6W���N�Cٺ��������� h�ҩ�!�`�(i3@��( ���M/*�3҇	��*��O`�� \)
�:qEp���,��\[��l�,t���H[W?��	P �a��e�D.7�q���f�e�M?��y�!�`�(i3����&��r��졾�g�Y������y�!�`�(i3�߆�p�h�T���ӄ��!�qgy�`��vN*���k� �ԬQ���Kͽ<\��1tSjv�!�`�(i3�o�t����w�`L����Y� �أY_���!�`�(i3i�Q�������=��w)��
=b~*��s�������P�íN=]a��o���H�RtV�^!�`�(i3�<@���ل=����h��'�j
/��ݚ�Н��Ra])n#���r����!�`�(i3�<@���ل=����h�Wsp[��X��=@'ѥ�
�:qEp�;�P�t�5!�`�(i3���F��O�VA�ڦ�c4
L	�\k]�x������ݚ�Н�
̛�]���n���G΂��b+}y[!�`�(i3]���\�x8���D�kJe���N�ScM?��y�!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3��jVѭ@!�`�(i3,�˳�*C[��l�,t���H[W?��	P �a��e�D.7�q���f�e�&�U��f�!�`�(i3����&��r��졾�g�Y������y�!�`�(i3�߆�p�h�T���ӄ��!�qg[���**���k� �ԬQ����5��t�1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=b~*��s�������P�íN=]8k��.ͥ�H�RtV�^!�`�(i3�<@���ل=����h�]
���7Ϝ�}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��OEʨ�`N/������&G!�`�(i3�7����������EN.74/�������yr�!�`�(i3�����!�`�(i3�7����������EN.74/���g!�%=F�=!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	������6��V(pyL0DMlE'�! !�`�(i3�<@���ل=����h�Wsp[��X��=@'ѥ�M`�K)��v�:�-22�v�I����~u/��kOT����1��eǡ��=֔׹���& d��]�?��\fʧ��sx�L<��}�u�?�d���&��R����\R��T;jZ@��2�c�n��`��O�W]�J#;?�k`���aF<��[��CC��z>9�R��$1&O^	QW�Q!r~$�}>���/�k�2�������P��d��1X���W߯{�����p�;����0,uD�*'�*of���вh��N�M�0��F{�r��졾�g��[��o}�����<@���ل=����h��g�:�B��K49�ݚ�Н�!�`�(i3ҷ��.G��-򅤅Җ��_j����EjP� �5ǖ�o�D���k$ !�`�(i3{�d"���ƍ2���lĸpAy����TRViY�ڥ����Ⱦ�<@���ل=����h��,�F��P��jVѭ@!�`�(i3!�`�(i3��b+}y[Z����r����%6��ڥ����Ⱦ�<@���ل=����h��J�m�X��-򅤅Җ��_j��� �ilچ=��X� 2!�`�(i3jꪑ��{�K�~�2��
 JSV`t�j�O��[��o}���P'M���k$ !�`�(i3?Q�@X>#�N-Y&yo�q΃/��}�y6�T�@�����M6�o8:4�g�G��0\��.5.\֯���,T���k�[��l�,���h<��K��I/����B�!�`�(i3!�`�(i3!�`�(i3!�`�(i3������P0�����K��I/N#~8"�Z��
��ܨCK�5uoЫ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3����C=+f2�s%���F��G�6{u��F�z�>�/� �=��Q�d�G}%����3f�B7�Q�+ż٧��jd�C���U�
{�~j9}^p�t|�7Ԝ7(u�!�`�(i3@��]V8ml�i��- �!�`�(i3�B�+2��;�P�ƺ'���g�;�jmT�#������PX6و�cµ L#_/�e��-����!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3T�=qއ*|X6و�cµ��%��(����e_�������B
�:qEp'{w#/ B!�`�(i3]���\�x8�:
1���Ư����z��>!XM�#����+1�;�.��1�>!XM�#�=5.B�����'����u��r��!�`�(i3h5���=�t���_j������'�.�Hh:��!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i3UI����������=��w)��
=b~*��s�������P�íN=]b~*��s�������P�ڎC�?�a%��w�ݚ�Н���+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ�!�`�(i3i�:`�+PN#~8"�Z��q�����8���&�
�:qEp'{w#/ B!�`�(i3h5���=�t���_j���M}����B�q�$x=��!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �m�ڨ�hծ�ݓ�W���q��n-���3��Y$��� л�g�G��0�-a0a3����|e"M`�K)��v�:�-22�vn��뾦��ݚ�Н����g!h!����e_�g�+C��sG��Hb� h�ҩι�+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ��q�9�ͭ�Ƀ�?PA�g�+C��sc�'�3<
���D�kJ��}Dq�f��߆�p�h�T���ӄM*QfY�"Z�Va�ir�K��I/��0�|�_�mS8<�n�ݚ�Н��7����������EN.�r6���`������ݚ�Н�ђw�)�WA�qIp��K/�k�2�]�u��y!�`�(i3��i��:q����J�sy�V��R�f+v�k�@duP���2�Q:��?��b~*��s�������P�íN=]I/��\]� h�ҩι�+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ��q�9�ͭ�Ƀ�?PA�g�+C��sU_GD��W�ݚ�Н���w�w:�!�`�(i3��Aڬ&W럼�~=�L�.ama�`m�5s�FF'l/7w|]/(繸P:$�O����K��I/��0�|섃Va�ir�K��I/z�
1���;G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��A~����>������!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEp���,��\���ևA�d��-��!��EJ��7o�*H��& ��0>!XM�#����+1�;�.��1�>!XM�#�[��l�,t���H[W?M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�a�݌3)�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�M���yt7�o�*H��& ��0>!XM�#����+1��*Hx�g�>!XM�#�[��l�,t���H[W?�>Jj:&ֲ!�`�(i3�A!���iW3��O�����%����:�������7�|���޵.��g�d�H�RtV�^!�`�(i3�<@���ل=����h�s��m�Eq�e>%����!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEp��`�ҪJ�F�z�>�/�a�'�Zy.
�@�����K��I/z�
1���;}2��L�)6g����O�Q:��?��I�^$D���������P�꠼*d�m����xQ�1tSjv�!�`�(i3�o�t����w�`L�&�����~��~\�Ԙx Ȇ�r��
!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�M���yt7�o�*H��& ��0>!XM�#����ևA1F#�֞qduP���2
�M����d��-��!duP���2�:
1���Ư����z���B� �b��!�`�(i3�7����������EN.�r6���`������ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sm@����K�ݚ�Н��Ra])n#���r����!�`�(i3�<@���ل=����h����3��[<�m��I�!�`�(i3T�=qއ*|X6و�cµd���2��C��C&��!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f�
L	�\k]ǩ�/f�]�!�`�(i3NQw
[��K���!n��뾦�!�`�(i3�U�Z^�t� "���
w�����z!�`�(i3]���\�x8���D�kJe���N�ScM?��y�!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3:)!�1%�@�	^���yCw�Hm���K��I/y�b�G2!�`�(i3i�Q���'���>;#��Z<��A!>!XM�#����+1�;�.��1���-����!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3T�=qއ*|X6و�cµ���(A�,"��C&��՝� s�#W���wL�'l/7w|]/(繸P:$�O����K��I/03�� <I��:����iW3��OEʨ�`N/�x{^4��*m!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3:)!�1%�@�	^���yCw�Hm����x�a�t!�`�(i31���~!�`�(i3@v��e��]�Լ�c���J�������n�0R��#���n��*ȑs>!XM�#����+1�;�.��1�>!XM�#�[��l�,t���H[W?[�G���K��4	_������=�#����=��'����u��r��!�`�(i3h5���=�t���_j������'�.�Hh:��!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i3��\7�f��T�g��� z�P��۶&��L�H��>E-�N�&Cd�c��aj�\iW3��OEʨ�`N/���:�������7�|���޵.��_�mS8<�n�ݚ�Н���+�t2��Lq��QF[�Z9�+	�ӸK)~� �ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#~x]V�{���>E-�N�&Cd�c��aj�\iW3��O�����%���	��$��\���@�<���7�|���޵.��N��:��!�`�(i3Yf����ڛ�e�D.7�q���f�e���	P �a�����=��w)��
=I/��\]� h�ҩ�!�`�(i3@��( ���M/*�3�IX�B��7����[j!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i36�B��~ ��A�Y�
���3ʩ�V$=�b�������P�꠼*d�m����xQ��q�d`��8]�Լ�c���J����
%�6W����!�qg�X�R&cE���-����!�`�(i3�D�������{
B��e�g��'�B�oSU!�`�(i3!�`�(i3!�`�(i3�T0�10#��vR�j�!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3��i��:q����J�sy�V��RkB�����X
%�6W��b�3�怜gVdxQ,�K��I/��0�|섃Va�ir�K��I/z�
1���;�����u��r��!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3:)!�1%�@�	^���yCw�Hm���\-{���!�`�(i3�����!�`�(i3�7����������EN.�r6���`������ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sU_GD��W�ݚ�Н�fĉ>99��A0ok��
�:qEp:䩒=]'!�`�(i3��:���r2Z�i��/79�O��F����{L,8�7�}ퟐž_�F��H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z�z��B��������p�:��q�՝� s�#���k$ ����l��T���ӄ��!�qgy�`��vN*���k� �ԬQ����5��t�*���k� �q� P�G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��A~����>������!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEpm���n�iW3��OEʨ�`N/���:����J0i�,�LD�s�x�-����!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>1�Ѯ�a�!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[�Z9�+	Ҳ�}�%Dܭ��}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3z�b۶p�t@�&|!�`�(i3���4)c�ݘ<�̆xƍ2���l�;�jmT�#������PX6و�cµ L#_/�e��-����!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3T�=qއ*|X6و�cµ��%��(����e_�������B
�:qEp'{w#/ B!�`�(i3]���\�x8�:
1���Ư����z��>!XM�#����+1�;�.��1�>!XM�#�=5.B�����'����u��r��!�`�(i3h5���=�t���_j������'�.�Hh:��!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i3UI����������=��w)��
=b~*��s�������P�íN=]b~*��s�������P�ڎC�?�a%��w�ݚ�Н���+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ�!�`�(i3i�:`�+PN#~8"�Z��q�����8���&�
�:qEp'{w#/ B!�`�(i3h5���=�t���_j���M}����B�q�$x=��!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �(*�O�qe��0�U������K���%>�rG�4���n�HN��R���IX0F�M��Eg�뚵]k�WM��q.��:�P9d^\'@�A2wKaC�IX0F�MV�ҁGG�K�BN
\�O.C�U��B��-F�}�WP'�uKwm�����"sS<GYqcHTX�';��#j�ݚ�Н��'�c��dN�<@Iv��nt=:��:5A��p~�vE�sy����D�� �v��}Dq�f��Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н��r$ɓ����˃�IG��Hb� h�ҩ������ya�E�Rq���my$�N��o�/���;
�:qEp'{w#/ B;�jmT�#�^N�!���<Ԍj��_�mS8<�n�ݚ�Н���\9"�ͱz�4��9m$����ˇ��:����
�ݚ�Н��,�3U�gN�k������ˇ��<��#�!�`�(i3��$F@S�� 63����1�m�
�:qEp'{w#/ B�&d,4���H��̣��+#�x"��g����0`$f��_Ub�F�S�1 �Бc�8-��E��B�1������}������!�`�(i3uD�*'�c�gyB��I��`j!�`�(i3��w�w:�!�`�(i3��.J7h�lr�{��|e��0�U+�qbp@�!�`�(i3HN��R��bP�63Z�t!�`�(i3�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�af��pD�Ё��
O�� ��A�Y�j<�i|n��$F@S� � ��>Bw�R���y+1�����8|��Rz�C�@;1r�S�ML�?l�Λ�~��o�fy�U��)���Y;e�iK-pm!9�>��n4s1�U��B��-��^�uJ#��r$ɓǉ�.y�U=������&G�7������JcH�����}�%Dܭ!��"� +}04~B3��������h��`�����y_�mS8<�nx��7��̖UB�no 2�X�h~������EN.��k�{����Ě���aT��3G�IX0F�M`�M�����> X2-�g����1���1X��94��f"����t�T��?E-h���U���e��_	�Ƽ��S�J\7 ��>�:�xjzӝ���w3��׍�&�U��f�����&���/N���74/����G🕾{�߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&G�7����׌�yt��\�k	䶙%;�������w�`L��t���Q�5ߧE4��Fr��jrc^Y�G�1X��94��f"��^R9��"�7�l5�5��U	�`�o��_�Rv�䩲$����E)e|A��`���φ��<�6��7�癆cgR������������ h�ҩ�i�:`�+P��=�ڹ&J�A7�伩���@|��璓�c�������t �[l;M?��yв��M$��2�w������vP8�J�g�*����3���E�i�m}6O�D mWN��ܐ�}������#�Ƀ�?PA �[k���?�Ƀ�?PAD��d�꺹_TR�\+�[\ٿ�6�P�`2����]'\gWg��	�Z�kfcj��r���iI9�o«IX0F�M�ȏ֦�"�\���F�`y������T�8k��.ͥ�Pi�#��Rk��H�"<�������$�\%e��}Dq�f��K��I/z�
1���;%��v�ک���&��m���d���ZMB���b+}y[^	QW�Q!r�TmY>��'�-��h��ƍ2���l�����C=+f3�{~��u�"ª���!��"� +}0�ʂ�j�Ï��	�l�lM�3 Pi�#��Rk��H�"<������ ��U�_:��}Dq�f��K��I/z�
1���;c�'�3<
�:
1���ƥ���W��D������0q�#�׾ŞWsuzS�n�(�a�ȠȎ�8��F��=5.B����Cw�Hm���K��I/@�k�F��ws� ��<C}���{��%��(�T�g���,�Ջ ��C�;�P�t�5�׹�3��܌o�l��������6�!&kݺ&m��
&+��[N'G�+R���o��_�Rv�䩲$��8��I�:Fa�7������A���!���;oN�	mH��7�癆cgQw�c4~Nr_�mS8<�n������ݰM�_�G]�;o�� ����nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r���_��*��j9�Y܉���a��o���H�RtV�^����C=+fI�#�ǖ����%��(��U�,��/�[9o������Ě����E�i�m}6O�D mWN��ܐ�}��B7�Q�����A@�yk�		������PsIT%�:α��2�N�3���!�qg��r�U���K���!q����`U�m���d�����W�B��C8�4�X�-}?�+������P�8�>�}��0�����f�r�wb3�@gò���S���"��gL
˙{�ʖCd��O|��������y���*We{4�ϋ�G)?2��H\�{4���I�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�ܸ�r��%W��*���u�Z�LQ[��Y��
�m��_��I�u���=���-m�N�cU���?*�����u��Ј�q%r&H�?�tUuf�ȖuB��x��=m��s׬k)[QH�x��E��_/<�_ ֻ��n,ꑮ'�J~72�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcdM�MQ l������W��ߜD��k�pqi��0	�J?,���Vr���F�!��c��Ď��J�c��[�R��0���h��\�ڰ�ȧ�`�>R�; i�V�JD�IX0F�MV�ҁGG%4vkz����`���φ��<�6�](ùy�;ShT���A(�c���_G��Hb�S����
̛�]��v�7b�%��v�ڕd�tu�z���?T��'�PD�����g�Z��3��a���!@�f")u��r��)Յ�N��I~F2�~H�c}��q_*�`�	a�F�������R:k�ڛ1���`��xm��s�Ū���l��A�k�C�!ax��]�z�[��CC��#\npu��r��d�tu�z���?T](ùy�;�T�TN��!�`�(i31���~!�`�(i3](ùy�;K� |�>�
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�^�#�nw�#�C����h�99^���+| �"R� ��ߌ�U��)���Y;e�iK!���d.d�G}%����3fU��KA��E)/�R��!�M���K�'ž1�|�'�����j��c�Q�n62�}�����\�X%��v�ڹ�+�t2�4\%��t����{�fR��}��k+Q�h'�Ȝx�5W ��̫(�H��
J��-|��Y��VF�˷��d��-��!g��J�s��F�e{iʖ.� �9�!��-������+�t2���<��������{���}Dq�f�E����[�k�n�=���b+}y[����l��A�k�C����.��y�� h�ҩ�`��v
K<�Y�|�8'�^�����ݚ�Н���Ě�����}Dq�f�-��)'�	�;���x��"u�����`�����>��-/a8!�`�(i3�1!�J�G�W�^�|�����NM������%>�rGO�D mWNfĉ>99��A0ok����Ě���P��U@Dφ��<�6�^���+| ���J�فN-Y&yo�q����,�ǰ	M,��rER�����Wݬ����W��P�Rn��EU���'���e{���Iv�z���AZ���d���!i^���+| �"��D�!�I�؉P-7i�J١����D)9W ֒���\�`��w9��x�i8B23`���x{�$��'!�(�JZ�Vk�;��|B[�x��ޗg�AOn�u?�!�`�(i3!�`�(i3!�`�(i3���aR�����Nh�NvpB(����揱�.FV�x�i8B23`���x{?Za����oA&��>���p[4$Ckj��������y��ܬS-l�ݫ&�b%%�Jם����2�wXw��<����f%T�^�c����L�{��:|O/�Ax�i8B23`���x{�CyW�f�tR�wX���V���G�8J��P>��t}�F��<�3y��������g�J�g�*�;^F�#�8 �X�G�[o�`��ۅ�e�\���Iz~r�;-�+�uM���X�\�{�4��֥��h>�p�c^���u�C^�Lc�V/��ﬄ;�%Ag�][ɓ4p�MRާ5a&���m��	6��L�W�]��'��v�|ӢBmi�>�/��z0�9"�{G;,^ ����E`6���3'�o�`��ۅ�9FhN�.�q��;��ƺ�3"�Z��ۑ�J��P>�TOi��;g��Cj��/	ol'3�Q��n�
ҍm�Euk�[�� �`�{x�<[�UXp�ߡ�?���	��V�j��S�n�(�a��kH���/֯���,&�7ݽ)g�G��0>߰�e��A�0q�#�ci߄��tw�t���_	�Ƽ��S�J\7rc^Y�G�K����-��h�r%��W���dB�Ro�F�tw�t����`UNP�_��1{Y�NY�]�2��ݚ�Н�#l'U:�g[/���^͒֯���,+�O���e���!
��g�G��0��p!�g>��ݚ�Н��K�,ǆ�`�܋�n焞 L#_/�e�!*��*8��!�qgg�f�p~(��|�x@S�n�(�a4N�J�ף������&G!�`�(i3U�07�:�tMɶ���74/����Y�G���֗*��ڡ�4-Y���Ra])n#����,��=7�7K�P�l[�Ƶ�	���QC�Ҷ����Sn	ͷg�?��R��3��m���d�0/0`9N1��-����!�`�(i3�,�B���{
Biۧ˺�s�˭;{o�Ϧ����ھ	!�`�(i3	���A��m���d�e���N�Scx��w����֯���,-}���A�I�^$D��Ҫ�\���S)`u0�F��a_�mS8<�n�ݚ�Н��o�t��8c���L���f�\%�+�8EN9��Z��.�\��$���w�w:�!�`�(i3��3�Z�#aȮ۔��5��Y��x�1�-Ϩ�ݚ�Н����F��O�/�"�����y?�?L�����������T�3��Y$�
̛�]��q00���龸b+}y[;�jmT�#��\���S)G�6�!~�������� h�ҩΖ7������8R ���M/*�3���\��/.f1]�?���	��x��ݚ�Н��o�t��8c���L���f�\%�+�8E��`�78>�٪�o�_&�
�:qEp�;�P�t�5ʁ���MյF:Ȱ����N9��Z��w���v��D�H����g�G��0��'���C&8k��.ͥ�H�RtV�^�D�����0	�+G�c��=����h� 8�2�~S�e>%����M`�K)��v�R�<<�U!�`�(i3'�^�����ݚ�Н���jVѭ@!�`�(i3�,�B���{
Biۧ˺�s�˭;{o�Ϧ����ھ	!�`�(i3)Յ�N���^�v�����;q��b+}y[���%>�rGO�D mWNG�&ց�*�&��j������ț}�	76�&�|��3��׹���& d��(�"x6�if�z�U��6T�k���#�;G�R��Nr�jfC��$�rˊv�����*ȑs;��|B<&ǒ8��#���H
�S��z��p2�������r'f�H��م���R7�j�2>����?XW�~a���@=�y�z�:���br� e8�~����d�4� ��@�1�˓I��#��pG|t�L7�="|k�{�:2��,���C� ���Б�����ph�)��ݯǖ���d�4� ��@�1�˓�C=�"C�@pG|t�L7��o��o����Z��O.C��>�w�Y�#E�m ��?Z��G.�w�ϸ��#|S������3[�u8�2W�+�?"J�L�Y\ٿ�6�PC��uB&ǣ©��A��4�h���6X�Obq0�~����O�΃S���ݚ�Н�*��^�"~Hv�"�ӏ$0Q���s�(�;�g�&�0m'�$p���=�t����}�(�
4��c��^�
E����d���m l�o�&�C�/w�x�P���E�`JcU!�`�(i3XO����0¤լq��/&M���<�q��9wS7��_�_��Kp�h�x0�7l]�) !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�0�����n!�`�(i3Y�"O���j����I~!�`�(i3��*�{6�.�ۊ䱃��ݚ�Н�.ӗ�r�(Z+�,�~�7!�`�(i3k S���zǣ©��
.�Ūz�/>�"�Ax!�`�(i3��3�N;C�]�'!�`�(i3��5@~Ju*k`Ë��!�`�(i3��)�ߜG���p�Gg,Z�fg�g���rz�!X�I�Y(��.�����R�!�`�(i3r� ��i�(���B��������d��$J�!�`�(i3%+bn/�{�.��8z�f������<��N�Lf�?ǉ�=���S���_�������"�9(���ԫrI�C�i�4��v�
 ��4���>�*�!�`�(i3���K�7��"hQ`� <�6�Q=)?`��BH2l}�{rcKE#���.�)�p�������s��+qѭ�+g[�</Sn��-�¾L��S��I����yP2Ni�~�ݚ�Н�X+&wG��	�X;p`�l.�	�C˹�+�t2��ӱ}�tMTl�����)��.��f�?ǉ�=<9����-����b=�`
 ֢��-�¾L��S��I���fÓ����ݚ�Н���퇇М1�X;p`�B��C8�4`�Z�l{�*������Э~���VczZ��������[�D���~�ߗ���@Tvs��&8�,��	�ݟȌ�V����f���w���4Wt#���'��(��8���/�f�?ǉ�=]a%ڔ�-����B@����u���M=�*������R���e�D�
�~��\��f��E��Ⱦʤ �� #��� !�`�(i3czZ�����ݫ&�b%%ׇӭ���1:	��?-����6��8Ͱ�����/���i� ��+��FI~u�#�$IXB2!n!����p
v�	�G���	(��7��F�dHG[��gR ��5/�`g��p&2P��KY+��1���~!�`�(i3!�`�(i3!�`�(i3?Q�@X>#�����
hxV��	��yϨ�ܛ9�~'0l�L�����}Dq�f�!�`�(i3!�`�(i3!�`�(i3��r�5�ѝ��泃�e{Q_�dbzL����ہ���M�!��^��BcƍItJm�Ԗ�Б�����ph�)ɪk^�P� e8�~��n,[������l��?F��٢�^���B0S�������*0]y� e8�~��*<!�F��66����~�"���D�tj�ڌMtY���l��2���:A�^���B0S �80D� �;��|B���r����!�`�(i3!�`�(i3�mJ�0�6�d=��¾ȼދ�Y"�I�,��u�C���L�s�ޘR�7h�,b0V�u�Q�ݚ�Н�b��
ߎ� n2ϒ�ȡ�&Y��V��G8T�w�nf�?ǉ�=�e�MW������L���	)��\R�][[�!�`�(i3�#�l+��B@
��B��+ H��*�{6��=��?��P�Y�6��!=.�
kZ)� [��v���Q:�7-mł(��gR� �ұf�?ǉ�=�;�.A�ى1�#��d_!�`�(i3�a\;V@|ऩ�jU/�\���WO+�jqh&Σ�h��I�
C���m�o��vPD��<!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�xsˁ�#2\z���L�f�\c`���6	D��&8�,�e'M�)�p��dHj�m�!�`�(i3m3�țZ��_�`I� B�!�`�(i3�<��N�Lf�?ǉ�=�$�V��bst�N���!�`�(i3�#ŪS�������k+#2\z��}�� �с�!�`�(i3�&8�,�e*���	�A�XF�����?UT>��˳����:=,3�/�r^�h!O���!�`�(i3frw��?�̞��>��vbëdP��_Ӯ\8�����$	�_:iO�A��*/�|��&8�,�H*W��u�a�ݚ�Н��>�@�C5]�꼧5#b|���Mk S���zǣ©���u��4��#�N�X�!�`�(i3�M�����{��A�Wu����������zq�{���r#�9l$H�RtV�^�k�O�>�dv��oTN֢&@��&�� ���)�{� �"�$�~c/kx��D(ކ�'T���+�ӱ}�tM�U젩`#�4>?� �1�z�����M�_~�:N���X)�:����s'-!�`�(i3եa�����苇��Fe#OOJd֯� ly����)�{� �"�$�~c/)R��L-���wӨj]h�u.$���8�$��`��Z���]�}��Px���A��4�h8�����ey�E���x�ր�ݚ�Н�E�%�� ��X;p`�����G9L�M�7��<�n~�<�&��Xh�hk��z���a��1�M]�!�`�(i3�G����/ӳxW8�8J�|9-B�U!���A��4�h���!U�020�$�~c/�*���J= �P���R�^=^���3�&8�,�6.���͈��?d��H���ź��*�3���g���/ӳx^Xp�ђ��ݚ�Н��֠������"���l<o�;)�y�y������x�������U/�e��<��(���B���A�� ��XI��/^�=O�gL뫵Ӷ�%�TE����k$ !�`�(i3!�`�(i3!�`�(i3��\a���_�x�BVo6;��|Bh�ƺ��y��D�m��
!�`�(i3!�`�(i3!�`�(i3�mJ�0�6�w�R���y��0�J���C!v���&!��U���0�+jq�����Å��������l=�w�����5�O�%E#P�$��Xo�Cn�g1�䁛����$�b9���dIvp@�J�y��*?(�oy=R.
�{� &�'�+�a8,�g�&�0mɬc��WN�鈑�)݁S�/dݪ�D�/?2�,ëYf�1�%A?�dL"� r�������7�����q�©�����[����YO�.Ŝϸ��#|S������3[�u8�GLa���mdЧ^{�j-����h��t���oޯ!�`�(i3��I�Ūe�E7.�Z�"�4��%�;��7���ө�Rxem_�$n����������������i�^�=���p��R�f�?ǉ�=�w�Ylj;!k�2Nc��Nn%{�oꠓόz#�<���X�u��
)\Y��!�`�(i3
)c?�%Q/�}| �e����kn4@Q�/��ݚ�Н����S�|J�X;p`�B��C8�4`�Z�l{?V��j�c�[N�&ѐczZ�����ݫ&�b%%f�?ǉ�=��=m緒6����}F��(ja]p�X�o|30��^?8�$��`���	(��7��P�v	��Y�Q9���ۗ&8�,�cop ���6�G|�</Sn��-�¾L��S��I����yP2Ni�~�ݚ�Н�*��^�"~H��
�[�<�`A��_i¼\K��
�:qEp0���Y$�8�$��`��7dh�?f�?ǉ�=�*46;�[-��$ϙRl�bu�	?�cx�3Lv	̅��!�`�(i3>N0Θ��ݚ�Н�Gظ0�����X;p`�l.�	�C�
�:qEp�����%������r��	��
�Q�}��"���l<o�;)�y�y������x���m[3�� ��
m}:[�O9UNTnF�\F�l9Z��b�Bϱ�\��FHѽ����8H���&�bP����|�J�=��?R�����!hh����P.���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3��kw�G��.�g3Zꢯ�wv��ޟ��}tt��wN�p%
-bK��:z6�U���e����T�bC�9/���U��)���Y;e�iK-pm!9�>��n4s1�U��B��-_S���\���&�vf��G���"sS<GYqcHTX�';��#jx��7��� �ؼ��"ª���!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^g�G��0��}�m�'�M �cJ$���hpI�_�c�r%�[�ap�Vȓ�"����Y�5ߧE4��Fr��j�p���"k��yV�:���(�'���:?���