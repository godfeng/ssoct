��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:�� �c�=0N���6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,xh'�$k�w�D1���}����ň���x�w�Y��k��ı���$��������j��t�w )�1��kN<��;��� B]�pE���	x]̃Dj#^Da����M�ٲ��9ߪ�
�M��ļz����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��Sd,�ϱ����@N1�w�0XL��t:w�~�gm��+��9��kT!����Y�f��a�Z��V2 �Q[6�i��<&�̝n�U��Y�C���t�#K�{ʓ��d��?�A\���5���a["<7U�i�#6u�,Уd�^:$�$���?#�+jN�N�{M}@���x�h�v[�2)ݛk�}dXQ������K����{Z�/*0�(bѮƷ��,�&'��Y_�68m}C��Z1)fd�vĻ�E����F5���Xf/���Jm�WH)5�Z!{����
F�P?_�!B�]M"Aw��-��ׇӭ��!�`�(i3!�`�(i3u0��L<q�`�c&�r.�?cXE;�i~p��M��gCu(o?C�����5	�)kJ#��t�{ڼ�`a3� �x���f:3���/�ky3�����=��ׇӭ��!�`�(i3!�`�(i3*8�2�z�����b/?�8I.���^r�b(�c�?����4����o���������i���%��S��!����P�><1N��r'�)d
�u|�$�iah7��f2`�r��sȸ�"rR!�`�(i3!�`�(i3R����G�ތ_tO~��E@�͔��Ġ�L �*�2R�W�~�26��\K�y؄@�!�`�(i3!�`�(i3/��oi�#��+��:iR��Sp㨚��}��6�8�-Zy?X��?��W���;��B�lXK�y؄@�!�`�(i3!�`�(i3�Կ���pu&a�vU0��p�$;�n ��j�ּ���)`4Zp��/���ϲ���>h�c}����>I	���(��B�:����@���4W�-c8��"3���s��ׇӭ��!�`�(i3!�`�(i30R��=	�@����W��nl@O4茸z���q����R��C���CS�� ��!�`�(i3!�`�(i3�0�9&،EB����n��|1�b�YL��&\VI`,xJ�����g}����&�������!�`�(i3!�`�(i3�>=���#9����'*�J�.�����G����%�,b�_�Ќ��*��4.���Xt�.U���ͧ�uQ0�})�����,]�x	��gf���{�P�1|5я����j���ֵ��sȸ�"rR!�`�(i3!�`�(i3_|?k��\+X��Y��8�-Zy?X�!�ZN9���2�䦒ccnh?�!�`�(i3!�`�(i3��j0��x���jz�H�gf���~�c��"��&\VI`, �DO'�L!�`�(i3!�`�(i3����N���z�����6u=�{��ZMN��>�! ,��e�w�1V�N��:˽�_k[9��~��!�`�(i3!�`�(i3'�Z�8�'��ѯh��d�J�\���=��&\VI`,f���a�9e47�O��C��_���U�`�R�Z-��شУ�X��d�rW��y����Fz�!�`�(i3!�`�(i3q<m6p��*u�j}@�El����WtUr���dp�
�2 ��Q=ߎ�����,������ccnh?���&\VI`,�=JK�t�J%�r �14�X#�Mwn5�����z1�z�F���ϡe����W*�RYS�Kh�!�`�(i3!�`�(i3!�`�(i3�q��L�!?�d���&�u&a�v��� a�ik��Wʍ3�V�޷��i�mm	�>!�`�(i3!�`�(i3!�`�(i3�@��ÂbݩJ�\���=��&\VI`,门:<#B�����+C���~KM�gzu4��	�!�`�(i3!�`�(i3!�`�(i3�U��a��*��>i�!i�X!�!D��(J�f�)�s�%�hH�oe��C��c�S+d�J�Г��f�u�����!-��B<ԧ�[��+��sȸ�"rR!�`�(i3!�`�(i3p{���gM�k���lh�&ĵ�	ƹqE_���RQ�
�)T^�b�k�@����S��l��ׇӭ��!�`�(i3!�`�(i3J�Y,�~)�{lN}Q�b�o�m��}�؝�TVq�|`kK��I�t����ۀ ��m��5ѧ��Z>)E�d��Z�����d�*���Fz�!�`�(i3!�`�(i3������!���C�/�y���ܴ�WM�P[��j�$�*7I���y�L�=sȸ�"rR!�`�(i3!�`�(i3+���6>�2'5�sZw��Q����}2M�; ����������-N��]�1�l0�)�Myիnň��h����]ߺ�`@��h�h����M����CN�u!�`�(i3!�`�(i3!�`�(i3��_�����v�����������U��5�D�v�l�Ū�TD���wG",���˫�i�m|� ��>K�U��L��nc�^��ns)��E�$�S��Z(�j�!wS����G�N�����ڭ�[��
A�4ϦE�6����ѹ��6[��{ֱ@����G��Mr�J�Mۀ7���\� ��2Rn�k�*��� ^ȣ�2$6�sI4$2�¤}@|��d��\��'ٽ$Id`ȯ~���Uz���+ߜ)��ns)��E�$d??�A��?U��|�����X�4V�.�(A���C�/�yV<��ϚEP�@�z���c>�I ��bv.�]0�[X�b\g!"�a$��z�e&Y��WM�P[��=����Vq�|`kK��I�`\�L',�y�+(̇�0S&",f�e��sƲ����e:ɄP���'㦡���0�8*��#�N�J���}��R���j�y���i�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������ݧu7Y�M�+|�#��Byl}Vİ�8�d��N��Ԫ^��rL�t��^�:AԪ^��rL�g�j�m��}��w�G���RJ��p�99-#` ������b_]s��2��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcfe./��:�!9\��N5�w��J��Zo  �0WP�da����'Q�:��~�z7	9��sE���ye��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#�.�x^ok��u4�� L�ʿԪ^��rL�Nl�Dvg�	Ԫ^��rL�t��^�:AԪ^��rL�>���x�<Ԫ^��rL�%�7��Ŀ<Ԫ^��rL���7�C)"�Ԫ^��rL���	��D9�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcQ#�y�&(���B��|/~.)��3\�R�F*}�c}��uO�^VM,q���\��K[�J�#��9�ĒTC��0���M�<lbtsR�b�"oʭ��4>rS��w�>��S���Fl�p�7Z0D@X�,4�?nϦE�6���������;%J���v�_�Q[�1��*��!?9�~����p>{��`�'�X�څ�˺�ƒLX���!I/���r&��\���%-��]�O���.e��!��z����)P����(��jD!���5�Nn>��
�*�EB���a�i #�� ��&��*mm�!=�y����h�}y(;⟝*#>*��4DA�,#��e�o?�M��;]��,��K!�ۻ2�e�1�ΟÈ�bH\�a�����RL�a)r��fI����F�����o�E���^�½w�>��S�Y�)\��B���|��S��2�)�Ln|����O2qs��s�L�:�;�T?��{}��+�����v�ɢ/*0�(b�ԝ���ɨVu��7���	x]̷?��+*�7��Mv�9�I��P2g-W~���џ�_�v%䨉͞N	����V���
��G'�۰�����M�,А�r냸�~���c�6�fST�jf&�~�7���}~�N{`1Kqn���D���i����	x]�)�RV!�7��Mv�9�I��P2g`X�8�\џ�_�v%䨉͞N	����V���
��G'�۰�����M�,А�r냸�~���c�6�fST�jf&�~�7���}~�N{`1Kqn���D���i����	x]���Ec��$7��Mv�9b�L-���MƝb*��4�8�:r&@��j�2Mk�(�VU)��*��u3����r���B��jN���7�� ��߼
�d�8DJ� ��m�!=�y����h�}jh�6g���_�-ִ�fY��/��Sd,�ϱ��Hx�U����� B�&"�D���i����	x]�����O��}�$L�7��`6�^���g&����a������}���D�"t�G�8=e����wHmM>p��&k��������Ԗ��RL�a)3���ʉ����H7��jX�+[�d�vԌz��S!�zg�Z�$e0���0��B�cN���	F�o�=�e �m�X������+�ct�ǈQ���\�4�s��{��]Q�TT	q��$��<�z5��J��eb�hW!'!7U�i�#!����P�>;�Ղ��G}Z��2�p��Oi�v���j�������JM�7")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t�	g�y�mq;����z��r���]��7ď%W�����k��d��&e�_�#�gWr���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QLi/-�#�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��'p�@�I�?g�f���\X�<����8��UWJ��)��q鋴�*Х�]��:K�E�\��Y�e hI�ˋ��vE-,b����Ǘ�Yзq8�Ј$�F5k0B�v�Ys�S�)�I,�D�y:d`A� ���8�TP���14�:v~E�)d,�vd���xi�X!�!D��(J�f�'��q�S<IÙ=�H%v@����f�7>�����ǚr��y��[7�d|���XP��ȅ&��3J��\G�Y#�u�'�'�7��r�=�����5	���]���>����C��U���e��E����Fv�Z��P,Nό���.ӻ���j��+`VU�2���HF3���̰�!w���B}�����
L'���Xw��E�d����N�DNl�@No��u��]�!����M[��Ǣ�K�&�a�*�p���@IE�U��>��l%i�-�%t̓�@��=�O��TD��ό���.Ӂ��̰�!_���RQ�
�����
L'���Xw�j�7���I,�D�y:#9�]�B��`6�����������s���,0=]^	�&|#9��Ė�{�!�`�(i3��(�
t�������2%=dϖ�i�q㧵�0������0��D��L���_�L�3��0I}.�?u����4�GO�L2�W�K����Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$:v��`E�EYZ/�h�@�o��I�?g�f���\X�<����8��UWJ��)��q鋴�*Х�]��:K�E�\��Yh}Nw���H�p0����1�, �>1�Pq�@\w��0]b!��u�=�?��3���Z�����]�!����w�Հ�(.V�����b��Mޡ.pz�Lۘq���U���g�,P�nw�����A�?���0yV�6IWJE�!r}<ﷹ�t�Z�f����@1��?�T�\ �ͻIb����rs�i�/ �m^'��D24N<I8����\.W^�V]��}R�wX��}�
�?�套�qD0t
�X��)�Bh����YW��b'�3AirW&IQ`�9�h@Zd\a�U4�1i�7�cL���	Ǹ�y85��6�S��y��Q{�^9�� ��¾�7܌:��0z�cUL��)���2N��n�O�3bg�������5	�3C���_����$�Qu������*�pf���rs�i�/ �m^'��D24N<I8����\.WPW���[f|#9����$�Qu�g��-����Q]� _�rs�i�@|`y
���T�\ �͜����Ƀd�#��Ӏ�`,9�H�Wa(􆿳��W��{q3�RD���Ɯ���:=��={���u�b�?9rscX{�X!,�x�������H�BnR�j�/T�<�_�{_8�Y��=�}�Vݨ��}Dq�f��x����մ�JH��j�/T�<�_�����fH�ݚ�Н���C�����Z���{�u1H3��)�.����!�`�(i3e )9���������$t���b�E�(�R��6�����6�o��D�muշ!Rq4���V�WR��4ŵݓ�W�����'%Ő^	ݠ�m��/N+0�-zNv�x���b�ʁ���Mյ���K,W�L?��:����
�T�z�D�RG�&ց�*�Wl�@���h�6�q��_������8���&�(*�O�q�
�+f ���2N�3u����V�*7��}Dq�f��x�����E!Ƙ�	�j�/T�<�_hv�a��Ww�ݚ�Н�{?�sce���Z���{�u1H3�^���3.�!�`�(i3��?���jA��������$t���o��/�3��6��D�Z��]+�D�mu�#��bE���V�WR��4ŵݓ�W���0|�.�ݠ�m��/���%��ō�x���b�ʁ���Mյ����
}�L?��:'��<X�T�z�D�RG�&ց�*憜��D�h�6�q����}j�4�8�8���&�(*�O�qe��0�U��2N�3u�sQ%�K�	��}Dq�f���4�CD5���}Dq�f�����M�3�@ym�2q�H�ﾅ1੡�3҃Cʅ��$	���z�B=�B���d]�B�H�� h�ҩ�P�d�=/;����-=B��*��O�t���	������$o���!�`�(i3!�`�(i3!�`�(i3u��>������\�S|��R[Y`8h��(�B��ұ��E���!�`�(i3".���X	"X�AUu���2a� 뻻%�qzB��W�w�\۹$I_e�8���/���}Dq�f�1���~֭�h��O=�bً����ȋ�H���RA<,�l�}�L@t�>��k��$f��_Ub��7��G_��Ct�w#��@������37y����m�/
?aT��3G���"��y�:����D<��5�2ԗ0z�cUL@Nr����d
z����YUr�(��z�jE��>��G������g�[�~���������g���^=�?��3��J��R���=�?��3�5�%1dg�(R\֎u��xp�"�/�(R\֎u�eK�	�$V�|ag��6��j�V��v�@x�2��`,9�H�W�I,�D�y:#9�]�B���`�6#��V��&�J��:�����(R\֎u�M+P��˝Sz��E�4.@�7��y%%C�+߮��5˚2�<��B���}�&E���m"`�7#���Q�X�<a|��6j�"Hs#�{'��#✲�@��P�6�}�j�GS �q{d�����5�:�ဳ��R����*k���pثIX0F�MF�� J�ʯ�7I���VjԿvU!�`�(i3�3FV�J�3פ����t��}pshI��Tޅiy:Vy�a���$�Qu�)�˥D@���f70����E����F��K�J���N}�m��{��b>�8�k(Ue-��C�-r��|ڑM��6�ZQ ��b�FP&��̘էHr�#�ڊ<?@��,۽��ֱ�q��e�X�·�fp�����!�`�(i3jݭ�F���%,�������;���EWre�E��5��!�`�(i3���D	��U~�&w���^�B���u�܎���x�*aE�ֱ�q��W$���� ��K�ł���f70���x�]�V���Oo��[*������%čr�|��B����g����W5OL�U����I��O.C��7�癆cg�ɨ�lܤ\�v'�w򻄸J\$41tSjv�@{s,����)P<�ܓ�Y.��J���&_��=]�RCJ�����@�ĵm�|#HK���ɱ�������R�ό�ङ�N�!�`�(i3��7`��R�>�3 �Q�/��@����*��Sx��1SX� �uE9�+����Q�Y��F� �:���G�O���wbk�$����$���]�!������G�/��@���V��*J ʉ݋QOE���k����[�e�!�rs�i��:5A��p� ͷ�	�<KSˇ��~q�`�	6��.��J�޺��:p~	o����Ai Ͳw���T!�`�(i3����0��Gd�~{��	=��a�O�e�S��'���Xw
�T�r�5��� л���'��
,�3 l��/��@����*��Sx��4p��F?�J�8�7���}Dq�f��0\� ��+�(R\֎u��Gj7�uzE���k����[�e�!�rs�i�F��|�'�&љ�0�#��u��A��?����9�Kf��"�+�Z�*�G�v_�w\�Lq..ө���i4뱢�\`xS%���y��lD���|�D+��Z�!��/��@����*��Sx��4p��F?�J�8�7���}Dq�f��%t̓�@���ʳ�(�	=��a�O�e�S��'���Xw
�T�r�5��� л���'��
���i���.��J�޺��:p~	o����Ai Ͳw���T!�`�(i3=�?��3�W�^�|��E���k����[�e�!�rs�i��:5A��p� ͷ�	�cp#`�?�!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3=aUh������}�pd=!�`�(i3�NA7�%R�W"���z�X@*[�]���9qj�xm�N�e�{�W!�`�(i3����a�~9��tf��!�3$�J�5'!�`�(i3q�\E��0N�]|-������:Y�{'%sk����w�;{�'8{1�'��!�("|�7>�����ǚr��yݲ�Z��*�!�`�(i3����١�&X��!{}�IWA,�L�_���1tSjv�!�`�(i3�]��/ݐ�t)�9����K�ł��
�T�r�5�!�`�(i36�c���EN����"�q�l�J8C�Y�{'%s��F�6?��!�`�(i3EOJ�uxm�PQ%cp��g݈��,Ŵt�MyފVZ鎬�������(���%��@E�t�o��t!�`�(i3�k��^�1�]��g3������ɤ|c*�n9ie�{�W!�`�(i3����a�~9��tf��!e�E��5���:5A��p���y��lD�ۢ�z�*���e������w�w�vE�I�9�O��F�u�F8O*�E��J�����1��� �U��֜��3*A&-�Ri!�`�(i3x9�U��=�b�\=ï�-��4�1tSjv�!�`�(i3?V��j�c1����?��~l�d��)P<�ܓ�Y!�`�(i3�Ra])n#���r����!�`�(i3w�����A��ߎ�x��y�g�5��z�?D�8��!�`�(i3��Ě�����}Dq�f����%>�rG40�RS���$
�)!�`�(i31���~!�`�(i3���L2��500q~Ig~�կ	��@�u!��Z�G��8̀��P1��TmT9w�[:��q����%>�rGO�D mWN���%>�rG�E`���!�`�(i3�;b�-�2��;�P�t�5�Ra])n#���r������5j���"��ӌ�r��Ě���Ib��LI�#�vzR5�<5�q��e��u��r������*c�:�3���nu4Bޗ��;�fޟA'������s��R7��Owu�+Q�F �e�M'��Q� ~�����F��O�������
�1m�(�Q������ޝ���ð�&��0�`����ǆ| c�]h3�G�'�s2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcm���D�'!