��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�*���g S)�-E��N<��;���Z��4d��{�
��|��Ȋ)zo1���á�K���b��j.~���m��+���%	v3"C��dKBE7\F���r��C>C�݂�N$��/���	�0���'v6�o~�a�(E
PIU��>v��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&��t�7H��'jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��V�)��[�P��;�� 9�/�<"����_quf�tg����_��9(?��lds£����&��ix�AH�k[�^��_͎��T�k ���������	x]�<���eQ���X��\���|�@c���Կ�:�%n��e�ι̕��R)U�~�O���`Y�5���=�zX4P?�o��ľ��UW��͌Tfu��w)�S �J���vy7��Mv�9�h�s����b�z�Y8�:r&@�	��Ϸ)�����V\~{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�T�`�7?�\��4�/�I����D;�~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/�R����+��T��M��j@�����nEAНC��8��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hG[��{�ĘX�������_�~/�F߼
�dr���3/7D�d�/+M���"��ei,l����Fv!.�僢�#��i����S(�Z���kv
�u��7+�����I�>g���#�W�w��fD�5����`K�P�C�s�&R�߷�C�Q���clׇ��I�����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�!�hM�-�kǾ:op�n�j{	�	�%!�
c:�/� �����\����Y@�P��c�C����E���&�N@�q�#~.���\�爱�vL�vO�ډ�g���?i����k��u�� ���$���&�F*���o����"��C�\�ҬO�'�/��(�g
��������=�G�w�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�AJ�㗲F̞��>�F3�v��e	ʆ�In��tw�?�b�>�ʆ�In��t����s�c��B��r�� ���t�����kE�����B��!�>��y�3əLܒ��i����2��R���R�BK���Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �_d�Jq/W��]���mn�j{	�	�%!�
c:�/� �����\����Y@�P��c�C���w�xDp:��I�^�5��+8{�7�D�`����)��o|��S��u2�_���`�?�b�����[A?H��Z�!
���>X�J H��K�zk�����x<Ep�����BS��I�JT�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDLY�m��?H���la�|3k>�o|�?|(�Ԑ���e����޳[��g6�w��*��� �2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���Q���t���"��N��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Ј�q%�2���AIq�!������T]����΅�F�6?��߼
�d�3�tD��F3�v��e	�H`�ɕ�����a�"Z鎬�����}�f���� nqҺ�I�ju8xC���^!��\�z��J�@ N>�4�
���%�z_=����8H
k�F3�v��e	"���Zx(ޒ֙f���>cӯ�����{,џ�Ӆ�)�<1i��|:L:dK}g\���N�VjL*� � �����"��y��b�h��5க�p���q7�F ��`�k`3�M�lr?���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�Je�˜�Z�u|w��cv	��v���pKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��/lt�3�ʆ�In��t�\�Ȟ�S��T�V|;����"��y�L�*�g�;F3�v��e	�愉V﫞��fS���'K�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�IK���+�F��4��*۫�<����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�g�E���IA�Z�6�"K9��k��p!���?cC��O�-w��^l���Q�>4�b����"��y�0u�9�J{=�
�o���d�٣��c�A�L'~�8�y<b��������>��l%i�-���"��y�0u�9�J{=�
�o��xZ��j�
�a����c��������jƓ�[g�E���IA�WG���ڽjZk�~����p�l$���96v_ ��)�,T*O����開-�J4p'�>��\��:��Z鎬�������(���w�?�b�>��]�!���٥���E�c���w?�����XR�[R*$�s�,�TMo������a�"Z鎬�����}�f���Z�!
���m�]$���~����p��+��W��5��<�>�┈�����"��y��!���~�Z27B>q��T��h��<�q�P}��O���D�RD;���;*��I
�M&wZ��8y�D��ӎ���Pw-�h���&��t�F߼
�d�\�5`��3�Z27B>q��T��h��<�q�P}��O���D�RD;���;*��IɬcMē�����l���5�Y�w����9�<���N>�4�
����(�.P�3XRt%3�o2C�g�kgw�"��I66�v��Gߕ�bȃ�J�&[d���玣b\r�r�7N>�4�
��F��iW[�`����C}���D����q7�F �}x���c�є��E�tAO������D8�>V��ƞ�x%/���]���b�~��pj6DU}��S3<R�0�xZ��j�
�a����c�4t���d&Fo����W�3~p�����O�k���LC���أ�"4$X���2(wUF�|u�VUĻ�3���ne66�v��Gߕ�bȃ�J�߼
�dȱgW�48�\ wg���>��8�4���M��_(����@N��B�)Y�Pa�DQ�����BP�m��+���%	v3�u���k3�7DY��S�\6��L�͒1�:�Ω�*���g S)�-E���`&�`�y-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc؆-�qh��J<P���f�o'
���#�l�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I]�I�rT�8&\})����ai.���@��8���i�E̳&k����_/�A"�U���w�c*����N��N�.`�Z�����èV$ Hl�]���'�PD��R'cf���_ľFW[��(���Zj���
ŵ����n{��.�[�Ѡ� h�ҩ�p��xs�S�+���A�T�fĉ>99��A0ok�?�JY�)�Y`��jD4��S��c��څH�8��)8��~��(h(���B����Ph���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h9��)�N6��cN��������*�m����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�AJ�㗲F`�ю龀�k"Ty�,tT��A��蠿����d�Uf�揆0�бԧ2N��n���?���^��a�\����Nf[8��(&�L���p�`�6��Qu���% gWVbT+xΣ�}��Q?M8�f2���u�䯄���\�˺�KA2���ݚ�Н�
ҭ�3���]_�t?	�$f��_Ub��7��G_��Ct�w#��@��������"sS<xF��]@� h�ҩ�
ҭ�3���ߋ����-�;�P�t�5�37y�����:���b��qe� ���t�]/�b~�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����_c'�E�uv�8�����*�m����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開Ht7s��֨M��n������B��!�>��y�3əLܒ����D�i
��$�Qu�&�<��G�jݭ�F����μ<�e<�^��XzHL� ӃV5+��:��u�Y�KG�t4~?����:=�X��wB�ɬ�ݲæ����KA2���ݚ�Н�
ҭ�3���bo N��7����F��O�}�	76�&�R�Q���~��p���웂���a�"�_���3� �d��f~�	$�*]�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h����D]4�AV% h�|!�x��02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a/����N4Ҩ,Ű����!d�h��<�q��7܌:����3Eֱ�q������m�q�>1�Pq�@\w��0]���8-|�Dp��xs�S�3�Q=o_�}�w֒��S��c�ط�¶�`�aT��3G�#b"d�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�16P! ��"�{��K�n,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I7.���K���xc�1e><��B9�f�M�q��2!K���ž�N��� <&�M#<.�_&|"�ֱ�q������m�q�C��l"�u�$1yy_a(􆿳��$ڿ��Fյ[+8�-jI�etsb�d"L�X"u�UA.1tSjv���'T���+t�'jf�|sb�d"L�Ɯd� (�f퀔����`0�S�����N�|�("0�i��$��lq�0�+��J@�h�����XX�HN��R��bP�63Z�t�R'cf���R�\<۳�B���m��h��7�p� ���:=��1���h��&�R���f�+��}���E�i�m}640�RS���$
�)|�
h��sb�d"L���"X��[����fb�L�8ɵ�6�������ݸ����:������|�h�'��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcޒ*T K��(�W,�qlW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL[U�7�tW2�_%4Yȵ�ixUS�w�?�b�>ތ@�۰V��hC$?���;���EWr�AW˟������<�<���Ŝ��T�\ �͜����Ƀ�^��e��S�Ò�c�����u^,!Y�R�">_X�;P��ĆjS�O��b��֔3�lf,wKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�hBބkᄽ�K��d�r��N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開�/���VDq�`'���蠿����
���HK�0,���U<�d=��¾ȼʥ�nr]Y�$>�A�]�Q$i�~)A�aK�(zL�H+�4Э�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���){]O�d��oO+۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d;�"�7� ��5}�Y7s�9���o��S8��@糺뾃7܌:����3Eֱ�q������m�q�>1�Pq�@\w��0]���8-|�Dp��xs�S�״$(�>g���=�g���>��8��-�Ϡ���:=
ҭ�3����#F!�QO���w�_fHN��R��Gu�"�0�R�@�6�֐����o��4q�I�w�o���"��y�0u�9�J{=�
�o��xZ��j�
�a����c�������
C�4_�k�2N��n���?���^�7s�9���o>��l%i�-��èV$ Hl�]��"��ӌ�r7�%M����� +<�عU�.�;�#���Yk�����]]=w��S��0 ���(����W0�]��x@�������a�"�_���3�>�<�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��0/,ύ�@�|�2�v�r�G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y|�
�xr�ȳh�L>sP"G�wk��a�S.l"�S�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3���/��kOT�i7N�_	�z�w.{��w�_��(�6k�4d�{j��b�ڐ]���!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW���T�Ŭ��!^�̖g_�3���4�듴,`Y�{'%sa�6���� <&�M#'���Xw��`UNP� ��b�FP&���P��'���Xw�8&���I���|I�D�{�:���Qu���%��,�,
((�H*�iH��[��(��Ƹv��*Qx}�������m������E�i�m}6�E`���ʥ�nr]�b�N����LE�ZKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �EG�b�$;�!�%rf�c���;t>
�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڲ2ꧧ��*���xoϼZ'��io��@8w\�ĉ	��c''����:�ui���?8���yB-��fx���{�h�)ȗ�bB˶s.RO�#C�R_Ax�.��Cɹ��e�P�~V�t ��7[�ck�?4�V�ʄ�Z�^i�a2G�F���������\��:��AԢ�a\�w�?�b�>޼�\�v�	�+�&I(&�L��R'cf����T�x��QU���^4�;�jmT�#*m?mp'ǷG��Hb� h�ҩζ37y���#�&��S�#fĉ>99��A0ok�?�JY�)�֬w�J%�H�[�ӄqB�>�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������]�#0�f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vch��\��f�U���e[�.��<PM�Q�����-�s�<���dL�t+"r��T�M���v��]�#�Ϡs[�Vo	����j�K��&�|8�
a]���԰66��)?��B'm���4.���Ryt��'^�����������開A�]Y��[����kEP"G�wk��a�S.l"��<�W�C%��p��:յ[+8��i7N�_�Z9a��q����G��)ѳ��(�NT�|#HK��P�s)B�
u]9�#�I��-�����y��j��kr#��w �:5A��p���F��O�}�	76�&�R�V�"�0ɶ37y���}�:��4q�I�w�o2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����z���x?�q��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��B2�:c�G�&��T� �,��J�X�u��.tƎ�d��R��;���!oc�_W<��=�n��O���DƯu&7���F�!�_(����@҄���G��A"�U���'���_�)����u"��	�I]���d=��¾ȼuD�*'R�"0��<5�����}Y��	}�@��`-z����:N�:�לQ?M8�f2���u��o�t]`!�ð��T�ݚ�Н��r�@|�T�(چ���9%����M�$f��_Ub��7��G_��Ct�w#��@��S��c�ء#h�|4�q�T�4(����H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����{�'��1��}�Φ�F䘋N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開=$��X��a����xZ��j�
�a����c�4t���d�Zb.�Z����$�Qu�&�<��G�xZ��j�
�����0��X�I�����8-|�D��=�g���>��8��-�Ϡ���:=��1���h��&�R���f٫6�k��C6�Ϧ����u��A�0���򴶽!��\�Ж ���-3���B�1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�ϭ�Ϝ�f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX��DU}��S3<R�0�xZ��j�
�,(e�%�<��t��\��
=z�.(!�`�(i3!�`�(i3d�s��cqŸ��?��t��3D�I��5ֱ�q������m�q�P w�mz�����<RD§B ���`y�����n4s1Յ��:��~��,�,
((�H*�iH��[��(��o|���P�����Hk]��xR)Z��E�i�m}6�E`���ʥ�nr]�a�n�AaT��3GҴ�0�^�k�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcF�Z\�5w{�ѵ���1f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX���`����F���L�{�B���}$|~ïSup�xg쬉� }�ֱ�q������m�q�.4g$�co��=��ەI7յ[+8�Ǎ^�~��Ȓ�ߺ̆(1tSjv�p��xs�S�;�U#�s�RJ��#���jVѭ@Ƹv��*Qx?���P��%�E�i�m}6O�D mWNR�@�6�֐[�%�g�7O�j�M��2(wUF�|��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc[I�#M�n�����z���R��kBޫ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��Ʊ���0
r���h�țՇ_���ˡ�#��I��3���ne66�v��G���V>�R<�2N��n���?���^��b9���t�Kh�޴���clTn��.��|ȃ�+p�WHZ�a���2#�kH�RtV�^���]]=w��w`��q�Y$f��_Ub�G��VO�����3�}@��9�ڮW�S��?��L-�:��c
Ү��p7^��t�>��o�r� ��J��ݪ�j�޺�5%-�b�+�