��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�4��s�A�|Ԣ��g��B���������'Q�|FV;�SJ�)�Y¹w���j�Ѩ+_D)�}«^�Ԛ;Q����|�?]���p�����^��bg�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�fh>�F<}���U��d@��o�����\ �cG��Q�	}���bS�N1�	N�6��������t�
�-�M���w�1�l��=[���헧�d��r�6b��lY�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_��c�W_QL�V��늈K`��$�dR����.�D���J7"�?�0��&.bN�<�B>p\�?;�+C-\:HBm��+���V�^��T3���i�I�?g�fP���o7cWp��!5� �+8���K��_q'����8�b�^��\68Oy
��/~.)��3\�R�F*}�c}��uO�b�^��\'�	<Hmb����@k�ZV"���:��#tC���,?a��Q\�_qť��[�޿�Pb���ym��+�<4��ˌ�ň��h��֑�/6K�R^|p��� e�1�:�Ω�s8�R�	�}����pn�R��}\^�N����{jϾn]���
�C��n�%G�n|���S�BgVֶ)�tc��Pb���ym��+�ވΦ�籢ֺ�9b����@���Z&��i1�F�\��ۧ孡4�^|p��� e�1�:�Ω�.�&ʺr����$l2�W�K���n|���.r-����G�^|p��� e�1�:�Ω��#��,�K��ۭ�a;_�H�0$�r����;�(8h$�_֎��I�?g�f}�(g����n�Cac�J=�%��Gx$�r����;�(8*�wc���^�\��z�$�r����;�(8��p8�J���%��Gx$�r����;�(8���t��~�I�?g�f}�(g����6BOy�4�ǿt.C_����(Ҝ�qc��[b����@�W6r���["�=�bB��bg��B���S��I�?g�fP���o7cg~GW����d����=�� F:��+���!�`�(i3�i3<�f�D���X���`��wl��h��"u����E0qD�=�JHn��z���z�O҈;�$�?��(x+���1����@A��{�OF8Ј&29]��\G�YH�W�h���Q�#<4^��E����F��j��\w��0]��0�&�ͭ�h�O�0N�By3��<�]�!����M[��Ǣ2�����Vc2�����Vc�d���N)k� Ɓ����[;�W�@���TBd��pO�`�Wi&��]2�y�Z鎬����s(Ǳ��Qu����к?� fX!Ev�dB7@e��xG�I�d���e�ѵ�퇇М1!�`�(i3�����
L'���Xw�j�7���˷���T�\ ��:E��]��8֯���,ٝ5��&�]��-��%M-�`��8�4+0$�oI�K���;�Ӏ׌u�KI̊C��3EF!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�;�
Ҷ�R����!~�ĵ�.V!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=KO֔��S���k��]�yRy���4𢜋S�n�(�aO�LYw9���TD��-�`��8�4��3{�WW�����5B`�j����t�}^b
��<!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDB[i3[\iv�dB7@e�ݐ��ItP:x	wyE �2�w����~��iR�c7G#+�Ǘ0z�cUL�I��6���T�\ ��F6�Ʌ�ej�`^��M_�y�":-�Ϛ�aa�G��1Ǐ˨�g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�A���=���j�*y�`��/��D�|6�	}x����!��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3������#R�ᐐ��<ilYݙ�?��Ϙ`nd�d�`��S^J�Z�E����F7G#+��3L��'99�q�V'�M=���&������Ԕ�p!!v*!���OjV��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�沯ϕދf2^R���dv�
c����;覨��F�֒���\�!�`�(i3��(�
t�ژq���U�Y�4Eb����"-�&<`S?wh�6�!s}6,o�}a�C�Ǐ˨�g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�5#<Z�D���� aV��w<����=��8!��[:��'l:}��Q2�����Vc�@�Q�3�=�<���>k� Ɓ����[;�W�@�����C=+f?�a~[�B��]2�y�Z鎬����s(Ǳ��S�䡢��y��A_n�V��@�!6RRǬv!�`�(i3!�`�(i3!�`�(i3!�`�(i3H�,�]� ��:
1����$���qǩ��V���7E6�D�xW����C=+f�N�Cٺ��v�ј�"��Z鎬�������Ӊ*ݰM�_�G]���������-��%M�rs�i��s�٭��[Ø�;�x��`y�����V9{)=5.B����Y%T��BPe.��xu	�L$�����//��kOT������P��2Dg����|g�Y�'���Xw�����C���V9{)�����p������e.��xu	���S8�P?_������Cҷ��e�r�J�n���'�#&4�����7J�Ru?{��_H��lC�!�`�(i3!�`�(i3!�`�(i3!�`�(i3(z�>�Ր�Q��k֤�[�B�)���Ԕ�scX{�X!,!�`�(i3!�`�(i3!�`�(i3!�`�(i3R��:��IU�~�*�hz��W���᢯��0���%N
˚�W�T ��x���� �+��T��VM ���ރ��t��Lq��"�$"�N�p��G_/~.)��3<�鶰.��I��7�O���,��B	a"����몝j@_8g!�`�(i3����u��ʆ�In��tݯ
�WŁM�����~Z��_""�,�>E���	h��IB�Q�!��H�*.�PS���ۏO���qh����d,�;/�"���Z�>)����GAџV�T����g��L�*��l�|���j�tcmN���*��<����-[Z�N0[����	�v�]wɭ�7��r�=!�`�(i3��|g�Y�'���Xw�������펎��{5!�`�(i3c��Et��q���U��D�pc�2�����VcP�qoNK�s��}L�9k!�����^��g�u.$���!�`�(i3��|g�Y�'���Xwd�n]N٢R��F�D�g��U-�e�,���6+��c�r%�1�#��d_v�ј�"��Z鎬�������(���Wi��Ɔ�f ��*��mx��Z�n��[��{_8�Y��=�}�Vݨ��E�d��",oMG~�Յ$�O&�c��Et��q���U��*�p9��b�^��\��[|��w��T�mT\-!�`�(i3!�`�(i3!�`�(i3!�`�(i3%m�\�u��I�z�]NW���:j���Բv�+@!�`�(i3!�`�(i3!�`�(i3!�`�(i3D�k���?�8c�	�^�贅����	^����5���C��ЙMǿI?�ʪ%��1��(�
t�ژq���U��O�^Q��h���LDY�P|�gd#v�5�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=WlF��8�j�6G���8i�qcU������~�A�qIp��K7��h��;	��-��%M�rs�i���	�>�g��U-�e�,���6+�2�����Vc2�����Vcb{�o��Ш�G��g� ��^�5��^	QW�Q!r��$J�L�ԥJ	?a��j��\w��0]T#�3�["�",oMG~捕�tP��ؑ@IE�U��>��l%i�-��+g^l�h����M��"B��$I��w��,c�A�L'�{&j���O
�_�Z)|#9���T#�3�["����:� %Z�P�c@IE�U����S8�P䴰^MWܑt�h�Ҕ�1�L�+��8���/��.aX�bAKj�V��v��[H��p��(�
t��Y�{'%s2�ew�a(􆿳����^��x�j؀O��u`Ʒ%kYl���#�]�!����M[��Ǣ�\�2��s�6�>u�t�a�]2�y�Z鎬����y��|�!�p�uF� y ������J�2��b���w�x���� �+��T��VM �����:穞#S���D[�K����S��I�?g�f��R"N\����_�FD�ȝ�xE|!�9��V���|�'����Bi�p!�`�(i3��|g�Y�'���Xw��}Dq�f����ꀍ!�`�(i3��!%���ouD����ό���.ӏwbk�$���7Z��!�`�(i3c��Et��q���U�x��7��Z��M��
�	^���y�T<9 =��ui|Ɏ;�0z�cUL�I��6��7�C��zC@�:5A��p��\���S)| ���j�/�@TP3C^�㊉�	��q���U�x��7�֕iK�D�b=| ���j�T<9 =��ui|Ɏ;\w��0]�N��W���|	�WI!�`�(i3���
��3��]���>����C���0�&�ͭ�y{N�En�"�,�>E���7���Z鎬����7.~t=� ��U���e�!�`�(i3�Q����z��l�q���U�x��7��֯���, e���T'�ʓv��ui|Ɏ;\w��0]ݑ���&�d���%O�	^���y�z�ȃ�� ��]���c�A�L'@����g��'Uy\��x��7��|�;�Ojz���)e��'�ʓv��ui|Ɏ;\w��0]7�wtMM�ʪ%��1!�`�(i3�z�ȃ�� ��]���m^�=͹ǿ��W���ͽ�ʇTf�\kJ��� VU+I��vMb��s���r���x����y����D�,�H�JP��|���ْ5
�8��1�:�Ω�s8�R�	�}�����`h�ag������T�0��r2����u�UC٤(U���*#�!�`�(i3c��Et��q���U����?�@�|+l~�8!�`�(i3��|g�Y�'���Xw�����U�ЂDa��(���o�d�!�`�(i3��|g�Y�'���Xw��������P���Qi!�`�(i3v�ј�"��Z鎬�����	�7 �#Z��M��
�	^���yN�By3��<�]�!��	Ǹ�y85�����F�>R�wX���D������^́|�A!�`�(i3c��Et��q���U�[��N�������l�x�f7﹏��|g�Y�'���Xw��+x�r�2�6�d�f!�`�(i3v�ј�"��Z鎬�����X���*�����:(�L��%�U�Yl���#�]�!����M[��Ǣ[��l�,1B��CSk�"B��$I��w��,>����C��(R\֎u�J�g�*o3��Y߁t@IE�U����S8�bM� 2)G��8���/���E�d��",oMG~�Յ$�O&��]2�y�Z鎬�����	�7 �#��i|�l5R!�`�(i3Yl���#�]�!���D��L#���W���ͽ�ʇTf�\kJ��� VU+I��vMb��sw�Y��k��ı��*���q{?d']lj�޺�5%��m�+��
J��@���D��L���_�L�Ȳ�V�溜��D�,�H�9� I�,�-fce��,\ަ�It��;���:d#���>잣����i��E����F�'n�^0o�0��wU�g��Q������4��k�y'��a��u*K6H �i7�sp>g�?o�x^[��
Bq0�[X�b\g�##qYw�J��g�U�/Ax��R�>(�I��P�O���������G����<E�ªY0�Б����!�`�(i3"�,�>E��4];ˍH�,t����t�i�lK�軧:pPFy���U��!�`�(i3�E����F���8�TP���{��XT}u��Q��eF� $���v�]wɭ�7��r�=!�`�(i3N�By3��<�]�!����M[��Ǣ)�k�4�U!�`�(i3�����5	���]����,�JL����?D�8��R�����!�`�(i3�����5	���]���>����CΌh��eZ!�`�(i3Y%T��BPe.��xu	�>��l%i�-�5`z��s�Ƀ�?PA�':E����j���0z�cUL�I��6���T�\ ��:E��]��8S�n�(�a�x�f7﹏N�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�����5	���]���>����CηxmQ,ۘS!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FH=Y��@�E����F7G#+��\w��0]�o�t��F�e{iʖ.	��A���TD��ό���.Ӂ��̰�!i�q8�2t�ݡ��1����(�
t��Y�{'%s2�ew�a(􆿳����^���(R\֎u�,��7-�)�V�3j@IE�U��>��l%i�-�jo�'q�!�`�(i3�E����F7G#+��\w��0]EOJ�uxm�j��O" w�"�,�>E����-��%M�rs�i��;m��"xd#���>��CyW�f�tR�wX��q�\E��0�Y$�J��;!�`�(i3��(�
t��Y�{'%s^;$v�P��<�4�����6��	���`y���+Ќn'I�+��x�v/cs�x�f7﹏�����
L'���XwI<��f�E�#D�����Ә�N^��#;r�����S��I�?g�f���\X�<����8��U��Ĭ�һ��w'Q��u���k�ȻD�ou�*Y x�Sk�ZV"���:��#tC������s��Z����UV~s�"y����S�����5W/�؏�<
DN�"�,�>E��ʆ�In��t��Q�]��-P�vȜ�[��CC�n̈́�zL͊�q��]��B�����`��������6�Q��l0��F��j.��h��u>a�Ĝz�j2�4y������旔+�ez��2��2V��y �a�/�b�!�`�(i3!�`�(i3!�`�(i3!�`�(i3F<����x]}��q=c���U�>ŔBU��o�e�W�@c5����m\��FHѽ����8�b9���P9b��e<����g�M�v���r�E����F}�=Ll�����&}0�@nRFC#r��k�pqi�������:��H���o���&�t.�}g �N9����T�>��˳���:��N׾!���G�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�<԰4�8�0)�kE���[%Dz�a�!����[��C��"�,�>E��4];ˍH�,t����t�i�lK�軧:pPFy���U��"�,�>E��4];ˍH�6iQ����L?V{��\G�YH�W�h���Q�#<4^��E����F��j��\w��0]��0�&�ͭ�h�O�0N�By3��<�]�!����M[��Ǣ2�����Vc2�����Vc�d���N)k� Ɓ����[;�W�@��ϋ�LΗO!�`�(i3�]2�y�Z鎬�������(���Jם����"X��[��Q[R�7I����hoDy����L��if�icZ鎬����s(Ǳ��a����+���%GO�Y2*꧗|i�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3py�Ks2'���d�k��)�:�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���u �D����R��of��^��W�5܊i�;J���hB;��i|�l5R�]2�y�Z鎬����s(Ǳ�����O��*��Jyh����{0YafH�RtV�^!�`�(i3!�`�(i3!�`�(i3!�`�(i3*�m��Cl2���Gʔ,V�(f��r:]�k9i�:`�+P��[H��p�����
L'���Xwd�n]N�/��A���G�f�ȑ�)MyӚL��H�q������
G�a
y���m~�^�]��'!�`�(i3!�`�(i3!�`�(i3!�`�(i3��@dr�8�Ny�s�g�"��a=�P�?��ԭ�O��Un{�$�C��!�`�(i3!�`�(i3!�`�(i3!�`�(i3��R�ji4���k�

g�����k�WvO�$�ꃬ㽶q^���+| �g�YӅ:Ԭ����
L'���Xwm��5�������p����8ǒ�4ه�������{0Yaf��tA��]�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��$��Ґ�:���qʤ���-��Tz�+�E�Dtf���E����[�� �����Yl���#�]�!��3{ح���D��r'ىn����H��6{�$�˽�L��"k@:G�pP_��G*!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л���O)T�;e���p�����"��lmeI�Qj`���*1���s�lI2�����Vc�	�1�G�{qUte�\�������V9{)[��l�,���0Q�@IE�U��`�-9v���]�+贕>��E��yxN䙌�@)�d��a�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�Ɔ�X9�,��pZ�ìb!��u�zٺ��ID��V9{)���+1�=D��p7�e.��xu	�>��l%i�-����C=+f�B����>v�ј�"��Z鎬�������(���Jם����"X��[��Q[R�7����C=+f+�ýpv�ј�"��Z鎬����Ĺ#{���.aX�bAK�T�g�������_����j��<ͧ�:|��b+}y[����C=+f��>@Qթ�v�ј�"��Z鎬�������(���/��A���ތ%Ş�W�z��GQĪ/���=K��<_I!�`�(i3!�`�(i3!�`�(i3!�`�(i3%m�\�u��>��k3���^�����i��88Q�4��0:��r�Ů�!ev�mS��0�
���)�*Y x�Sk�ZV"���:��#tC������s��Z�����z���ْ5
�8��1�:�Ω�s8�R�	�}����pn�R��}L�Y�͋�<Ct�z&��â&�3ݾw�����$G⃍����,ԯ���gn��Ab�%^�;-оk�	ܷ�4D�Ps��܇�`5��\�vňu�,�s�?�/�2@V�����*�P�1ߒg�A�/�����%>%�����2 � ,w	����[7�d|���XP��� �vBX�y�E�e����KoϬ�ί��#�ڊ<?@��[	J��;I<��fҮ�w�Z�M�_F�k-�!�`�(i3�E����F��j��\w��0]��0�&�ͭ�h�O�0Y%T��BPe.��xu	�>��l%i�-Kp(����2�����VcƮ��.J� ���rqϟ<�^�5��q�\E��0!�`�(i3�E����F��j���0z�cUL�2�c�L��lC��U�T�\ ���A����u�#�$IXe���b���|g�Y�'���Xwd�n]N��F�dH����y���	ܷ�4D�P�r|�֖j��T�\ �͘�f��p�b�z'hۉ)��d�7�qĕ%t̓�@�H�\�{\�"�f'�gܜ�]���>����C����Wj4��⍽аN�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�]2�y�Z鎬����x�#w���Ƀ�?PA�c��|[��|g�Y�'���Xwd�n]N�/��A����Q[R�7Kp(����2�����Vc;��2h�����	�rl0�G�ņrŀ!0���!�I%H3�j�V��v�˩��*��c��Et��q���U���V9{)����0��G5���S)��TD��ό���.�^	QW�Q!r�#✲�@���K�*� �7G#+�Ǘ0z�cUL�2�c�L��lC��U�T�\ ��oR��m��%�э�g��L�*������
L'���Xwd�n]N��F�dH����y���	ܷ�4D�P�r|�֖j��T�\ ��oR��m��%�э�ghR�P�����
L'���Xwd�n]N�/��A����Q[R�7��+g^l���v�Z�"B��$I��w��,>����C�x�j؀O���ўC�k�Yl���#�]�!���D��L#���W���ͽ�ʇTf�\kJ��� VU+I��vMb��sw�Y��k��ı���$��������p侢���|�پ�`5���S��I�?g�f&:��r-,�/�����,��B	hI�ˋ������$G⃍��������u����\�vŽ�u��|Cݮ2����|�G�]R#�����ݱ���������u����\�vűhFyu�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�֚��IV�Tୌ�}��s�$����n|s�)>�vNd�)i!�`�(i3!�`�(i3!�`�(i3!�`�(i3�e/W���.�#���[�l�)��|B�;�h���}둮N�pS��Y�׈PzO�l>o��|�w��Y�ڪ!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDVW�ȏ�k��a�s+�ҟ�r/�^��D途��[��7�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=$L$E�͆صE�����&��Z�4���>��ru��!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=Zʓ�p�i�i��О	Q��J/[f�ͪ�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���w�>zɳ�B��,��C-2�^���ij�IRO�=���f.K!�`�(i3!�`�(i3!�`�(i3!�`�(i3�d���a�jwi�U���gh�䊉��	��J�6���G��"�WɆ&6�\]�4�6�t��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3؟��)�`U
]�,J��)v#��������6f1�W�`t��9��V�9!�`�(i3!�`�(i3!�`�(i3!�`�(i3WPtA��ro��� zv�۲=�k2gh�䊉�䞘gx�n�A��S� �WɆ&6�\]���x��MQ�(f��d;��,���O'��E��4�T}�Ĉ������=���f.K!�`�(i3!�`�(i3!�`�(i3!�`�(i3Ta�F�O���^�#��\�'L(\Ӧ�H�W�h���Q�#<4^�"�,�>E����-��%Mό���.���|��pe���b�Y%T��BPe.��xu	�>��l%i�-��9��稕!�`�(i3N�By3��<�]�!���TZ��Pj���$5�?� �٠Fd���e�ш�_(x��`!�`�(i3v�ј�"��Z鎬�������(���Jם����"X��[��Q[R�7D�wP�/�we���b�Yl���#�]�!��	Ǹ�y85��3}�@�7"j���b7xY�J��-4��h�]8e�0
A���J��@��^�}� u��=��5W_R�{ɟ=:�ْ5
�8��1�:�Ω�`��G��L�Y�͋�<Ct�z&��ÃlO ܅doGa�젿��ʐx�?WA{I�Z�T�����N\� n��A�T�g�v�;�K7���'n�^0o�)�?�^�?�XW������w
��ڎ:�ڛ)
�}��ɣ�YV�PD�E${��4`�˨�;O8�d�
~�n�}Y�:]�@�<g��ũ,+$\�M��lJY�Pt���`��8��f�`��[��Yt��'�d"[~6����aD6&>��Y��q��f�}��`<Y��sp�����5	���]���c�A�L'�������W��_�ړ8���/��4��}�<�N컽kg����|g�Y�'���Xw�j�7����'�e���"j���b7|#9���Y��
�iC�E����F��j��\w��0]%��C���+�
�c�~��j��\w��0]��0�&�ͭ�E����F��j��\w��0]{k�h�+m��q'��7G#+�Ǘ0z�cUL
 '&1���D���J��8���/�;9�".<�x���� �+��T���.��Б���뒴-UR�{ɟ=:�ْ5
�8��1�:�Ω�`��G�����R^| 4�,�-fce��,\ަ�Itnh'yt�;U��֜��3�:ET֤vKzL͊�q����ϡ����pܜ!�I�lW���LWɆ&6�\]j}8o{:�֕ߝԀ�I�R���F��c��Z��}��	�d�bzP#�-������4Q��#��w21�X��|�C#/<���q��!�u�ǭ��k��?��}��7Q�� +@��牥��*[���Μ���a�M+|�����\��6fz5�WRj�.(Wx*q�\E��0�v�4�oK���-��%M�rs�i��UQA$��5�%]���a(􆿳����^���2jɸ�����5	���]���c�A�L'�������W��_�ړ8���/�}T���y~:���_EH��o��C!T*�q���U����?�!�`�(i3c��Et��q���U��;���)"����}���c��Et��q���U�ЂDa��(o��0��7c��Et��q���U��ꢤ�Og�ШT�7V��(�
t��Y�{'%s���䒼�W& s��Ѩg��U-�eE������(e�0
A���J��@����S�BgV�0�ם�kj�޺�5%�ȻD�ou�*Y x�S���Z&��i1�F�\��ۧ孡4�Z�NCIw4t�iZ]XF����������'�e����ʺ�;[��\�v�W����ĮfA��x�%�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�GW���!��������F�┠�Gj���X��XM��d:p{�imlK:�� +@���0X�K�9D���o�j�0�J�vt�OF��������g2Uo�H�0�{�?Nt�!�ei�P�?��'&�s��Ia�|���+,�)��R�ᑧv0-�(4��AYpǞ��8sU��֜��3��TG���PIÙ=�H�c��Э|;>bv�E��5�F��������5	���]���c�A�L'�������W��_�ړ8���/��4��}�<�N컽kg����|g�Y�'���Xw�j�7����'�e���"j���b7|#9���Y��
�iC�E����F��j��\w��0]%��C���+�
�c�~��j��\w��0]��0�&�ͭ�E����F��j��\w��0]{k�h�+m��q'��7G#+�Ǘ0z�cUL
 '&1���D���J��8���/�;9�".<�x���� ��8[0p������arG�n�����KY�ʃ|�پ�`5���S��I�?g�f�SL�<.w[!�� Q鹈��fq�]�Xy8��;6aJVlO/����\{F˯�+)��ʺ�;[��\�v�W����ĮfA��x�%�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�GW���!�C�ד�c���O}a Օ�M� ���g):�.�k�ꂎ	�F�; ,@�� �^�4C3��xk޵ǋe����C����3�u�g̽2�-�l��S&�@ߧ�h�~�g��2߅_���c��`��Cm{w �<��>:Մ��F�9����'*#�b�B���m��d�7���A�f3��m��'A>�:ET֤vKzL͊�q���~�>2��p�ϵ�DEG�p�P�� nU�IÙ=�HF���m¡���r��1�Z���=���u*K6H�mV��5f��b�x#2���p5�}�]���x�]�V���KD:�}��lȻA��^8����̇i�d�?�c��Et��q���U����?�N�By3��<�]�!����M[��Ǣ����K? T��j��\w��0]KPkqy�{��
�%v]<��z��}�\w��0][�л���7��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<� ��i)Y�I��w��,c�A�L'J����l�!�Y�7#�xI��W��_�ړ8���/�;9�".<�x���� �+��T����)�G�o���sp%r�M$�*|�پ�`5���S��I�?g�f%��h,�qc��[]�Xy8��;6aJVlO/8֩]=$�G�p�P��g����="�,�>E��ʆ�In��t����Z����oY��8�b(��!�`�(i3Y%T��BP��&��J��bF���w¹��<d���<
DN�!�`�(i3�i3<�f�D���X���`��wl��h����f		d��2)�Yϰ0|]<w:�,ԯ���gn����fԱ@ι��QG�����U��!�`�(i3!�`�(i3x�]�V��;���Ӧ��Gjh�rO-�7(OK�� �"���
�v�u��̒m���A�/���a
%���A�+0�l�R<�jЉ/8y̚[b�0<���E����F��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+"�,�>E���TD���rs�i�jf� l�Ǜ������CyW�f�tR�wX��hs�����n��0�5	x��(�
t��Y�{'%s�:�f~=g(���B��ɓ�~Ҡ	u{ᵿ�����"X��[��Q[R�797*�SC�E����F7G#+�Ǘ0z�cULd�g>57<�b:m�X`�7���ө�)�F��3A�)Oqn�����ea�g��U-�eן�-�Q�Z�0V32;5�Y%T��BPe.��xu	�>��l%i�-|�秽m�E����F��j��\w��0]A��4�h���n�܀��TD��ό���.��l\�6�'����7Z���(�
t�ژq���U��s\���7�_~�:N���|g�Y�'���Xw�f�VHF��Q�#<4^�v�ј�"��Z鎬�����X���*�Lt�2�tN�By3��<�]�!����M[��Ǣ&��s���q�����5	���]����񁫴}2;9�".<�x���� �+��T��Rc1"�>_�q��.���{ᒺx�E'��:9�+�m��+^
s��mpM4,��=ٞO��q��f�}�����Hh�E����F�ҋX����>��l%i�-̇i�d�?�"�,�>E��<��z��}�\w��0]%��C���B��+ Hc��Et��q���U���5�G
mX��u22�7Ê7�E�4'���Xw�^�Ҍ�!�`�(i3N�By3��<Z鎬�������(����
Y�	�u*w�A��˦��<�/t�c��o��C!T*�q���U����v�� �!�`�(i37Ê7�E�4'���Xwd�n]N�7�����?�$����v���sY�ƹ@t�	��j��{l�f|�ό���.�4�3/Xδ!�`�(i3�����
L'���Xwd�n]N�7�����?�$����v�-��u��h;��!"�]��(�
t�������2�~�7���	��D܂�A�N�p��G_�(����5�6ԊM$x->J�"��Y����m�+��
J��@��sSL
��l�"�DUޑK��឴�����9����ۙ��\n�i�Z鎬�������(���2/
e�C�Yu*w�A�V9_=('��h�d �'���Xwd�n]N�W�R�ٶ�P �ZHA^�Xt��t-�]�Gڮ4\{Z鎬�������(���2/
e�C�Y�l�@qN=
��N�?�_u�
���)�*Y x�S$�r����;�(8�	S����x���� �+��T��#��=��v�����gT���Ai� �	{��E�D�|{�o��C!T*Y�{'%s2�ew����Tu��"U����I������L��{l�f|��rs�i�չ���m�g��U-�e�Æd�MS J�5�s��(�
t��Y�{'%s2�ew����Tu��"�I�r�?�q�1Ig� VU+I��vMb��s����v��9��zc�ds�gp�im����S��I�?g�f}�(g���̀:���o������L(\Ӧ�?�|����o��C!T*Y�{'%s2�ew����Tu��"U����I��Ly	I�"�,�>E���TD���rs�i�$ݝ��6�(�%�8����{�=�c-�����<YF`?7G#+����w�V�"-4��h�]8e�0
A���J��@��sSL
��l�"�DUޑKv�7I+jq��"�$"�N�p��G_�(����5�6ԊM$x->EN׹�TشP�ZyV �	{����aҗ�(�Q�#<4^�c��Et��q���U�ЂDa��(o��0��7v�ј�"��Z鎬����F�71�B�������%������5	���]���>����C���w��E����F��j���0z�cULm��.l��g��U-�e��,H/���,�)�x�P�1-6e.��xu	�>��l%i�-Ly	I�"�,�>E���TD���rs�i��g�M8X�(�%�8���(���^�;9�".<�x���� �+��T��#��=��v��>�"[�<�S�����m�+��
J��@��sSL
��l�"�DUޑK�7�������9��?)�$�M�ET�����'���Xwd�n]N�?���iv��$����v�/w1z��ӊ�����
L'���Xwd�n]N�W�R�ٶ��I�r�?�q�1Ig� VU+I��vMb��s����v����4W����ZI�6��ْ5
�8��1�:�Ω��#��,�GkO���������8����H���O5|�"�,�>E��<��z��}�\w��0]��0�&�ͭ!�`�(i3��{l�f|�ό���.��6[��u�V�<�nbBI��|g�Y�'���Xw�^�Ҍ�!�`�(i3N�By3��<Z鎬�������(����
Y�	�u*w�A��˦��<�/t�c��o��C!T*�q���U����v�� �!�`�(i37Ê7�E�4'���Xwd�n]N�7�����?�$����v���sY�ƹ@t�	��j��{l�f|�ό���.�4�3/Xδ!�`�(i3�����
L'���Xwd�n]N�7�����?�$����v�-��u��h;��!"�]��(�
t�������2�~�7���	��D܂�A�N�p��G_�(����5�6ԊM$x->�K�����܊ȻD�ou�*Y x�S��9����̠�P\�I1}Kط��4q�������o)�]rR��ӟ-���r�1���X���`��Fb��҆7���ө�q�#���Z�>)��<H�-��*����Kp&�@���k���a�\����9�	��%ι��QG�����U��зq8�Ј)w�<�_N���i��I<��fҾ��9�Ǧq��G8��=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A�����
�����Yl���#�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��kv޶Glbq�Z��T�I��w��,c�A�L'Qī�*pY��?� Zh�RG�p�PR��{�&�8���/�2�ZwŃ�9��|�����|g�Y�'���Xwp����B<�D-Ε�(�
t�ژq���U����?�"�,�>E����-��%Mό���.���|��p�}J�A��j��\w��0]%��C���]M��_�\"e.��xu	�*�QN����q�1Ig� VU+I��vMb��sw�mT� �j�޺�5%�ȻD�ou�*Y x�S�W6r���["�=�bB�K�E�\��Y�ea�;y� ����t���5���=\�B�wj$g�b9����$�n������ л�A�.�hQ3'�e�R��;�ݪ�򈟆�������\�vŽ�u��|E]�tM1-��E�}�?c7`��A�@c%��h�rs��l=�L)w�<�_N&�G"�2���k4I<��f�L(\Ӧ�H�W�h��e��|��j��\w��0]��0�&�ͭN�By3��<�]�!����M[��Ǣ&��s���qc��Et��q���U�!�`�(i3�v�d����7-ڍ�qL�\�b�`1���"3c���[���-��%M�rs�i��UQA$�R�^Ƒ����"X��[��Q[R�7D�wP�/�w�����	Z鎬�������(����U6�bL��W��_�ړ8���/�;9�".<�x���� �+��T����~��@�.��#=b��z���ْ5
�8��1�:�Ω�s8�R�	�}�����ֶ�#3��������K�E�\��Y�ea�;y� ����t�آ����<�bṪ�N��B�)Y�]V�H7'�U��֜��3JHn��z�ܐ{���E�q��f�}��h�'f R�E����F��j��\w��0]��0�&�ͭ!�`�(i3c��Et��q���U��>�w�Y�#���\��Fwv�ј�"��Z鎬�������(����F�dH�/�R�Ĳ4�������`y����>�w�Y�#+���G��v�ј�"��Z鎬�����	�7 �#�iK�D�b=4{W'M/��I��w��,>����C�pॻ}���E����F��j���0z�cULjaGkƊ~8����\.W^�V]��}R�wX�Ձ��̰�!w���B}�����
L'���Xw��E�d����N�DNl�@No��u��]�!����M[��Ǣ�K�&�a�*�p���@IE�U��>��l%i�-�%t̓�@��=�O��TD��ό���.Ӂ��̰�!_���RQ�
�����
L'���Xw�j�7����'�\�n`��!��B�T�\ ����NF��]� VU+I��vMb��sw�Y��k��ı����V���}����W*�׸-�nC/$q��"�$"�N�p��G_/~.)��3\�R�F*}�c}��uO�Go@3w��������]�Xy8��;6aJVlO/�4zG&/JD�*��z�l0��F��j-"{b���<#l=���E����F�_��������\{8����\.Wl0��F��j-"{b��]�0^ݵT"����S��i$ۇ��;q�:s�qDx=m��sEs��Wn2�B���s��[7�d|�Ҟ�%��bj�.(Wx*�_F�k-�!�`�(i3N�By3��<�]�!����M[��Ǣ���ꀍ"�,�>E����-��%Mό���.���C7}�7��r�=N�By3��<�]�!��	Ǹ�y85�B���0�1���U�<�o���8���/�-�}��d:�rQRтY%T��BPe.��xu	�>��l%i�-̣�^��!�`�(i3��|g�Y�'���Xw-�}��d�ܲ�k?Y%T��BPe.��xu	�>��l%i�-���!0%����Cs��|g�Y�'���Xw�P���w��:
1���Ƒ����E��@IE�U��>��l%i�-�%t̓�@��^́|�A��|g�Y�'���Xw-�}��dB<�L�V_Y%T��BPe.��xu	���S8�/ #O�)U��֜��3,0=]^	�&|#9����!\�'�ϝ�ˏiv�ј�"��Z鎬�����
��al>��`����E����F��j���0z�cUL���.�1�3�8���/�p����ݡ��1�������E��@IE�U����S8�P?_������`y�����������A�����"B��$I��w��,>����Cα��S&�r!�`�(i3��(�
t�ژq���U����������2Dg���"B��$I��w��,>����C��W�3�-c����L�{��(�
t��Y�{'%s��.|Z���ǚr��y�_��wBW��8���/���e��c<��/�a?�ґ����E��@IE�U����S8��<�J�QM����2�E~9���i�d�g��U-�e�,���6+��=v��� �	*�c9����"wg��=m��sD�}�*Uަ�_VS�䡼ڱa��NX��j$����f��׷9lD��XH�:ux����Yl���#�]�!����M[��Ǣn���H��5E^��Z�TD��ό���.ӷ9lD��XH:�b��t3Fj�a�k�]�!��	Ǹ�y85�������W����b~�>H7�v�ԯt*4�Z�"�	��D܂�A�N�p��G_/~.)��3\�R�F*}�c}��uO�Go@3w��������ǌL.��T��xdE���ƪ�M�D_���.���nEA��lRZ{%�