library verilog;
use verilog.vl_types.all;
entity altpll is
    generic(
        intended_device_family: string  := "Stratix";
        operation_mode  : string  := "NORMAL";
        pll_type        : string  := "AUTO";
        qualify_conf_done: string  := "OFF";
        compensate_clock: string  := "CLK0";
        scan_chain      : string  := "LONG";
        primary_clock   : string  := "inclk0";
        inclk0_input_frequency: integer := 1000;
        inclk1_input_frequency: integer := 0;
        gate_lock_signal: string  := "NO";
        gate_lock_counter: integer := 0;
        lock_high       : integer := 1;
        lock_low        : integer := 0;
        valid_lock_multiplier: integer := 1;
        invalid_lock_multiplier: integer := 5;
        switch_over_type: string  := "AUTO";
        switch_over_on_lossclk: string  := "OFF";
        switch_over_on_gated_lock: string  := "OFF";
        enable_switch_over_counter: string  := "OFF";
        switch_over_counter: integer := 0;
        feedback_source : string  := "EXTCLK0";
        bandwidth       : integer := 0;
        bandwidth_type  : string  := "UNUSED";
        lpm_hint        : string  := "UNUSED";
        spread_frequency: integer := 0;
        down_spread     : string  := "0.0";
        self_reset_on_gated_loss_lock: string  := "OFF";
        self_reset_on_loss_lock: string  := "OFF";
        lock_window_ui  : string  := "0.05";
        width_clock     : integer := 6;
        width_phasecounterselect: integer := 4;
        charge_pump_current_bits: integer := 9999;
        loop_filter_c_bits: integer := 9999;
        loop_filter_r_bits: integer := 9999;
        scan_chain_mif_file: string  := "UNUSED";
        simulation_type : string  := "functional";
        source_is_pll   : string  := "off";
        skip_vco        : string  := "off";
        clk9_multiply_by: integer := 1;
        clk8_multiply_by: integer := 1;
        clk7_multiply_by: integer := 1;
        clk6_multiply_by: integer := 1;
        clk5_multiply_by: integer := 1;
        clk4_multiply_by: integer := 1;
        clk3_multiply_by: integer := 1;
        clk2_multiply_by: integer := 1;
        clk1_multiply_by: integer := 1;
        clk0_multiply_by: integer := 1;
        clk9_divide_by  : integer := 1;
        clk8_divide_by  : integer := 1;
        clk7_divide_by  : integer := 1;
        clk6_divide_by  : integer := 1;
        clk5_divide_by  : integer := 1;
        clk4_divide_by  : integer := 1;
        clk3_divide_by  : integer := 1;
        clk2_divide_by  : integer := 1;
        clk1_divide_by  : integer := 1;
        clk0_divide_by  : integer := 1;
        clk9_phase_shift: string  := "0";
        clk8_phase_shift: string  := "0";
        clk7_phase_shift: string  := "0";
        clk6_phase_shift: string  := "0";
        clk5_phase_shift: string  := "0";
        clk4_phase_shift: string  := "0";
        clk3_phase_shift: string  := "0";
        clk2_phase_shift: string  := "0";
        clk1_phase_shift: string  := "0";
        clk0_phase_shift: string  := "0";
        clk5_time_delay : string  := "0";
        clk4_time_delay : string  := "0";
        clk3_time_delay : string  := "0";
        clk2_time_delay : string  := "0";
        clk1_time_delay : string  := "0";
        clk0_time_delay : string  := "0";
        clk9_duty_cycle : integer := 50;
        clk8_duty_cycle : integer := 50;
        clk7_duty_cycle : integer := 50;
        clk6_duty_cycle : integer := 50;
        clk5_duty_cycle : integer := 50;
        clk4_duty_cycle : integer := 50;
        clk3_duty_cycle : integer := 50;
        clk2_duty_cycle : integer := 50;
        clk1_duty_cycle : integer := 50;
        clk0_duty_cycle : integer := 50;
        clk9_use_even_counter_mode: string  := "OFF";
        clk8_use_even_counter_mode: string  := "OFF";
        clk7_use_even_counter_mode: string  := "OFF";
        clk6_use_even_counter_mode: string  := "OFF";
        clk5_use_even_counter_mode: string  := "OFF";
        clk4_use_even_counter_mode: string  := "OFF";
        clk3_use_even_counter_mode: string  := "OFF";
        clk2_use_even_counter_mode: string  := "OFF";
        clk1_use_even_counter_mode: string  := "OFF";
        clk0_use_even_counter_mode: string  := "OFF";
        clk9_use_even_counter_value: string  := "OFF";
        clk8_use_even_counter_value: string  := "OFF";
        clk7_use_even_counter_value: string  := "OFF";
        clk6_use_even_counter_value: string  := "OFF";
        clk5_use_even_counter_value: string  := "OFF";
        clk4_use_even_counter_value: string  := "OFF";
        clk3_use_even_counter_value: string  := "OFF";
        clk2_use_even_counter_value: string  := "OFF";
        clk1_use_even_counter_value: string  := "OFF";
        clk0_use_even_counter_value: string  := "OFF";
        clk2_output_frequency: integer := 0;
        clk1_output_frequency: integer := 0;
        clk0_output_frequency: integer := 0;
        extclk3_multiply_by: integer := 1;
        extclk2_multiply_by: integer := 1;
        extclk1_multiply_by: integer := 1;
        extclk0_multiply_by: integer := 1;
        extclk3_divide_by: integer := 1;
        extclk2_divide_by: integer := 1;
        extclk1_divide_by: integer := 1;
        extclk0_divide_by: integer := 1;
        extclk3_phase_shift: string  := "0";
        extclk2_phase_shift: string  := "0";
        extclk1_phase_shift: string  := "0";
        extclk0_phase_shift: string  := "0";
        extclk3_time_delay: string  := "0";
        extclk2_time_delay: string  := "0";
        extclk1_time_delay: string  := "0";
        extclk0_time_delay: string  := "0";
        extclk3_duty_cycle: integer := 50;
        extclk2_duty_cycle: integer := 50;
        extclk1_duty_cycle: integer := 50;
        extclk0_duty_cycle: integer := 50;
        vco_multiply_by : integer := 0;
        vco_divide_by   : integer := 0;
        sclkout0_phase_shift: string  := "0";
        sclkout1_phase_shift: string  := "0";
        dpa_multiply_by : integer := 0;
        dpa_divide_by   : integer := 0;
        dpa_divider     : integer := 0;
        vco_min         : integer := 0;
        vco_max         : integer := 0;
        vco_center      : integer := 0;
        pfd_min         : integer := 0;
        pfd_max         : integer := 0;
        m_initial       : integer := 1;
        m               : integer := 0;
        n               : integer := 1;
        m2              : integer := 1;
        n2              : integer := 1;
        ss              : integer := 0;
        l0_high         : integer := 1;
        l1_high         : integer := 1;
        g0_high         : integer := 1;
        g1_high         : integer := 1;
        g2_high         : integer := 1;
        g3_high         : integer := 1;
        e0_high         : integer := 1;
        e1_high         : integer := 1;
        e2_high         : integer := 1;
        e3_high         : integer := 1;
        l0_low          : integer := 1;
        l1_low          : integer := 1;
        g0_low          : integer := 1;
        g1_low          : integer := 1;
        g2_low          : integer := 1;
        g3_low          : integer := 1;
        e0_low          : integer := 1;
        e1_low          : integer := 1;
        e2_low          : integer := 1;
        e3_low          : integer := 1;
        l0_initial      : integer := 1;
        l1_initial      : integer := 1;
        g0_initial      : integer := 1;
        g1_initial      : integer := 1;
        g2_initial      : integer := 1;
        g3_initial      : integer := 1;
        e0_initial      : integer := 1;
        e1_initial      : integer := 1;
        e2_initial      : integer := 1;
        e3_initial      : integer := 1;
        l0_mode         : string  := "bypass";
        l1_mode         : string  := "bypass";
        g0_mode         : string  := "bypass";
        g1_mode         : string  := "bypass";
        g2_mode         : string  := "bypass";
        g3_mode         : string  := "bypass";
        e0_mode         : string  := "bypass";
        e1_mode         : string  := "bypass";
        e2_mode         : string  := "bypass";
        e3_mode         : string  := "bypass";
        l0_ph           : integer := 0;
        l1_ph           : integer := 0;
        g0_ph           : integer := 0;
        g1_ph           : integer := 0;
        g2_ph           : integer := 0;
        g3_ph           : integer := 0;
        e0_ph           : integer := 0;
        e1_ph           : integer := 0;
        e2_ph           : integer := 0;
        e3_ph           : integer := 0;
        m_ph            : integer := 0;
        l0_time_delay   : integer := 0;
        l1_time_delay   : integer := 0;
        g0_time_delay   : integer := 0;
        g1_time_delay   : integer := 0;
        g2_time_delay   : integer := 0;
        g3_time_delay   : integer := 0;
        e0_time_delay   : integer := 0;
        e1_time_delay   : integer := 0;
        e2_time_delay   : integer := 0;
        e3_time_delay   : integer := 0;
        m_time_delay    : integer := 0;
        n_time_delay    : integer := 0;
        extclk3_counter : string  := "e3";
        extclk2_counter : string  := "e2";
        extclk1_counter : string  := "e1";
        extclk0_counter : string  := "e0";
        clk9_counter    : string  := "c9";
        clk8_counter    : string  := "c8";
        clk7_counter    : string  := "c7";
        clk6_counter    : string  := "c6";
        clk5_counter    : string  := "l1";
        clk4_counter    : string  := "l0";
        clk3_counter    : string  := "g3";
        clk2_counter    : string  := "g2";
        clk1_counter    : string  := "g1";
        clk0_counter    : string  := "g0";
        enable0_counter : string  := "l0";
        enable1_counter : string  := "l0";
        charge_pump_current: integer := 2;
        loop_filter_r   : string  := "1.0";
        loop_filter_c   : integer := 5;
        vco_post_scale  : integer := 0;
        vco_frequency_control: string  := "AUTO";
        vco_phase_shift_step: integer := 0;
        lpm_type        : string  := "altpll";
        port_clkena0    : string  := "PORT_CONNECTIVITY";
        port_clkena1    : string  := "PORT_CONNECTIVITY";
        port_clkena2    : string  := "PORT_CONNECTIVITY";
        port_clkena3    : string  := "PORT_CONNECTIVITY";
        port_clkena4    : string  := "PORT_CONNECTIVITY";
        port_clkena5    : string  := "PORT_CONNECTIVITY";
        port_extclkena0 : string  := "PORT_CONNECTIVITY";
        port_extclkena1 : string  := "PORT_CONNECTIVITY";
        port_extclkena2 : string  := "PORT_CONNECTIVITY";
        port_extclkena3 : string  := "PORT_CONNECTIVITY";
        port_extclk0    : string  := "PORT_CONNECTIVITY";
        port_extclk1    : string  := "PORT_CONNECTIVITY";
        port_extclk2    : string  := "PORT_CONNECTIVITY";
        port_extclk3    : string  := "PORT_CONNECTIVITY";
        port_clk0       : string  := "PORT_CONNECTIVITY";
        port_clk1       : string  := "PORT_CONNECTIVITY";
        port_clk2       : string  := "PORT_CONNECTIVITY";
        port_clk3       : string  := "PORT_CONNECTIVITY";
        port_clk4       : string  := "PORT_CONNECTIVITY";
        port_clk5       : string  := "PORT_CONNECTIVITY";
        port_clk6       : string  := "PORT_CONNECTIVITY";
        port_clk7       : string  := "PORT_CONNECTIVITY";
        port_clk8       : string  := "PORT_CONNECTIVITY";
        port_clk9       : string  := "PORT_CONNECTIVITY";
        port_scandata   : string  := "PORT_CONNECTIVITY";
        port_scandataout: string  := "PORT_CONNECTIVITY";
        port_scandone   : string  := "PORT_CONNECTIVITY";
        port_sclkout1   : string  := "PORT_CONNECTIVITY";
        port_sclkout0   : string  := "PORT_CONNECTIVITY";
        port_clkbad0    : string  := "PORT_CONNECTIVITY";
        port_clkbad1    : string  := "PORT_CONNECTIVITY";
        port_activeclock: string  := "PORT_CONNECTIVITY";
        port_clkloss    : string  := "PORT_CONNECTIVITY";
        port_inclk1     : string  := "PORT_CONNECTIVITY";
        port_inclk0     : string  := "PORT_CONNECTIVITY";
        port_fbin       : string  := "PORT_CONNECTIVITY";
        port_fbout      : string  := "PORT_CONNECTIVITY";
        port_pllena     : string  := "PORT_CONNECTIVITY";
        port_clkswitch  : string  := "PORT_CONNECTIVITY";
        port_areset     : string  := "PORT_CONNECTIVITY";
        port_pfdena     : string  := "PORT_CONNECTIVITY";
        port_scanclk    : string  := "PORT_CONNECTIVITY";
        port_scanaclr   : string  := "PORT_CONNECTIVITY";
        port_scanread   : string  := "PORT_CONNECTIVITY";
        port_scanwrite  : string  := "PORT_CONNECTIVITY";
        port_enable0    : string  := "PORT_CONNECTIVITY";
        port_enable1    : string  := "PORT_CONNECTIVITY";
        port_locked     : string  := "PORT_CONNECTIVITY";
        port_configupdate: string  := "PORT_CONNECTIVITY";
        port_phasecounterselect: string  := "PORT_CONNECTIVITY";
        port_phasedone  : string  := "PORT_CONNECTIVITY";
        port_phasestep  : string  := "PORT_CONNECTIVITY";
        port_phaseupdown: string  := "PORT_CONNECTIVITY";
        port_vcooverrange: string  := "PORT_CONNECTIVITY";
        port_vcounderrange: string  := "PORT_CONNECTIVITY";
        port_scanclkena : string  := "PORT_CONNECTIVITY";
        using_fbmimicbidir_port: string  := "ON";
        c0_high         : integer := 1;
        c1_high         : integer := 1;
        c2_high         : integer := 1;
        c3_high         : integer := 1;
        c4_high         : integer := 1;
        c5_high         : integer := 1;
        c6_high         : integer := 1;
        c7_high         : integer := 1;
        c8_high         : integer := 1;
        c9_high         : integer := 1;
        c0_low          : integer := 1;
        c1_low          : integer := 1;
        c2_low          : integer := 1;
        c3_low          : integer := 1;
        c4_low          : integer := 1;
        c5_low          : integer := 1;
        c6_low          : integer := 1;
        c7_low          : integer := 1;
        c8_low          : integer := 1;
        c9_low          : integer := 1;
        c0_initial      : integer := 1;
        c1_initial      : integer := 1;
        c2_initial      : integer := 1;
        c3_initial      : integer := 1;
        c4_initial      : integer := 1;
        c5_initial      : integer := 1;
        c6_initial      : integer := 1;
        c7_initial      : integer := 1;
        c8_initial      : integer := 1;
        c9_initial      : integer := 1;
        c0_mode         : string  := "bypass";
        c1_mode         : string  := "bypass";
        c2_mode         : string  := "bypass";
        c3_mode         : string  := "bypass";
        c4_mode         : string  := "bypass";
        c5_mode         : string  := "bypass";
        c6_mode         : string  := "bypass";
        c7_mode         : string  := "bypass";
        c8_mode         : string  := "bypass";
        c9_mode         : string  := "bypass";
        c0_ph           : integer := 0;
        c1_ph           : integer := 0;
        c2_ph           : integer := 0;
        c3_ph           : integer := 0;
        c4_ph           : integer := 0;
        c5_ph           : integer := 0;
        c6_ph           : integer := 0;
        c7_ph           : integer := 0;
        c8_ph           : integer := 0;
        c9_ph           : integer := 0;
        c1_use_casc_in  : string  := "off";
        c2_use_casc_in  : string  := "off";
        c3_use_casc_in  : string  := "off";
        c4_use_casc_in  : string  := "off";
        c5_use_casc_in  : string  := "off";
        c6_use_casc_in  : string  := "off";
        c7_use_casc_in  : string  := "off";
        c8_use_casc_in  : string  := "off";
        c9_use_casc_in  : string  := "off";
        m_test_source   : integer := 5;
        c0_test_source  : integer := 5;
        c1_test_source  : integer := 5;
        c2_test_source  : integer := 5;
        c3_test_source  : integer := 5;
        c4_test_source  : integer := 5;
        c5_test_source  : integer := 5;
        c6_test_source  : integer := 5;
        c7_test_source  : integer := 5;
        c8_test_source  : integer := 5;
        c9_test_source  : integer := 5;
        sim_gate_lock_device_behavior: string  := "OFF"
    );
    port(
        inclk           : in     vl_logic_vector(1 downto 0);
        fbin            : in     vl_logic;
        pllena          : in     vl_logic;
        clkswitch       : in     vl_logic;
        areset          : in     vl_logic;
        pfdena          : in     vl_logic;
        clkena          : in     vl_logic_vector(5 downto 0);
        extclkena       : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanaclr        : in     vl_logic;
        scanclkena      : in     vl_logic;
        scanread        : in     vl_logic;
        scanwrite       : in     vl_logic;
        scandata        : in     vl_logic;
        phasecounterselect: in     vl_logic_vector;
        phaseupdown     : in     vl_logic;
        phasestep       : in     vl_logic;
        configupdate    : in     vl_logic;
        fbmimicbidir    : inout  vl_logic;
        clk             : out    vl_logic_vector;
        extclk          : out    vl_logic_vector(3 downto 0);
        clkbad          : out    vl_logic_vector(1 downto 0);
        enable0         : out    vl_logic;
        enable1         : out    vl_logic;
        activeclock     : out    vl_logic;
        clkloss         : out    vl_logic;
        locked          : out    vl_logic;
        scandataout     : out    vl_logic;
        scandone        : out    vl_logic;
        sclkout0        : out    vl_logic;
        sclkout1        : out    vl_logic;
        phasedone       : out    vl_logic;
        vcooverrange    : out    vl_logic;
        vcounderrange   : out    vl_logic;
        fbout           : out    vl_logic;
        fref            : out    vl_logic;
        icdrclk         : out    vl_logic
    );
end altpll;
