��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�S�T�;Ϗk[�^��_͎��T�k ������[���a�8%`��4�s�6�XAoeu��a@����þ�V�E`Ԏ��%��1��*�"��Yk"1/���%	v3"C��dKBE7\F���r��C>C�݂�N$��/���	�0���'v6�o~�a�(E
PIU��>v��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&���7�os!w����]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�K�MV}xj\�iW�(� 0�D�A~����p��ؚ�fD�~����pn��-�4ڭ	���
��M!�nz��m��+��$|��;D���J7"�K[�J�#��9�ĒTC��0���۞�^�� ����C��H$�ƵoB;sѱE�ouJ��p����B1�o3(�'�"̂����b4MI�-`7�(Y��;(��Цy���t��k�8���҆�|n�����|Hj`;U;�c=���)M�BJ�Й�m��/K5r��!����%�J l���&��RL�a)r��fI�����,�%��a����2��>҅eB���u���;��I�6r���ScB��\�~�q� \���T��U	�1�_u���V����*�^�~ì3"� �vm�!=�y����h�}��<]~8+|���g�S���!�<o?�M��;]l��j�z�	��A�b/���"��y�s����o�k�8���҆�|n����e��m*�~^T�ɴ�#���3J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|A�L�Y�͋�<��y�͌�4r�O��C��0��t�z�������_0ֲ�p����u���;�Թ!o�o,%H�%�ì���Tl�
� �AH���g���	]+��3�U�Z�a��w4hJ�=�ʝF@�4%�j�Fi,������00�m��I6�X'W�=������H�����/���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hl7�Fmi�E+���WY`�`��yZ鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QLi/-�#�
Ү��p7�I�?g�f�L#����2=�l����K�E�\��Y�9�{u��]�!��M8���	D%ϱN��ɐ�=%+]Bo�A;h�Fx��!��;�cY�~�ː<��cx�S���>��l%i�-<nvl*%ɬ�� ����y���+%:>п�p=	�˳͠m�xW�g]����n(���˧\w��0] B�A�wM��wb�S��V��^��\i�@^7&ģM�'n�^0o�<:�W�_�WzD9�G���:�����開�~������ZVG��т	�J�%�XB�&�=T-a�ؕJ�9�#=�8%T-a�ؕJ�>�5�0���6C�&/���_(����@N��B�)YN>�4�
��o�M���Z@0SDbz�@ʶ�橓[*jD�1Y�ΊS&}Z�F�>"�ѐw���5�W�u,�%UU��2��{i�X�x $}��}��uRBO ^�̒��b�|��@��l�
����gvS������H�|�ߦ��X�G[�Q��ǺΕ�Xw�} u�NT�<�*�!g()��ikp���H���JHn��z���}��-j�^�J��μ�\�v�w�?�b�>޼�\�vŌ�rf�Gѧt�� ���OgۈPM�����+u�VUĻ�3���ne��-���E�0w�m\+>���yg�E���IA���vsl�����p!���?cC��O�-w��^l���Q�>4�b����"��yvmH����{=�
�o���d�٣��c�A�L'~�8�y<b��������>��l%i�-���"��yvmH����{=�
�o��xZ��j�
�a����c��������u��u;xI|$�@(?udG���q�©���H��JnXe�+�Uz�QL���b{�"G�*ZkS0��N{a�9O��Yk"1/���%	v3L�Y�͋�<�B)�6��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�pv��[�\�)�A��m�aOLyb�7�a�`�2G%�/��Z>L}x��=��f0���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL���iM0�3y��#Q���Q�q��o
�X���C�~��~�Ln��S�W�ѐw���5u�0�yo�_���
.����Ď�rȫ�S ��Sup�xg쬉� }�ֱ�q������m�q�.4g$�co��=��ەI7յ[+8�Ǎ^�~�篯����hV$��-�����$�[��= -|�GP�ݚ�Н�
ҭ�3���#���1���b����@�Y~�`���Y-]�\^M�Ɣ�	��x��ݚ�Н�
ҭ�3���#���1���b����@�Y~�`���Y-]���v�9����Ě���!��"� +}���k$ ���n����-�����y��j��k\y[P޽��5 cd���%��E�/�xA���%0[-��&J��;b�-�2�'{w#/ BƸv��*Qx�!F�;^/K�2�+����e
,�p8�4��|r$J�-��^$f��_Ub��7��G_���;�P�t�5�37y�����:�3��s���EU1��?�}����0�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������P���2�z�I0���ԏc�r�(���7L��1�6`3bQ=�3��>�Dj�OgW���y�k�m2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y��� ����;*��k��J���\Ol����֑1Y�ΊS&�<�ɰ]�+��׌#��M'��P+V�_������o@i�1�P\�q[�7�����a�"e͉�Xk����0��hC$?���;���EWrf�Nd+l�Yҽ֗�1#��Z�����f���T,m����i�Ӛ��F�)[ Z|X��ٖ���g�OcH��9d���aX���$�Qu�&�<��G�!�`�(i37w|s���0�$i��kq?H^��2踫g(�r�N�ǁ�f�T��p_U
#yO�E���%�;���EWr�L�����!�`�(i3�b9���1]�?��� ��b�FP&��"��IJ�N�Q9�����-�)����=��ەI7յ[+8�Ǎ^�~�篯����hV$��-������"�=�X|�\dG��&(i�/B�\3���l�c1���~��DFTޱ}���0|Q�>8�ހ�$f��_Ub����b���잸��u��r��>���(���;*��k��� ��y���Y-]�[�Q0�M�1���~_'R�4���%�3�F�������78�4��|r?\�z?Xk�:䩒=]'5�����}Y��	}�@�r�<Uee�N������*��vbsQ?M8�f2ݜ�
N#�0���:s����"��IJ�N�Q9���2��n�v��/��@���#��M&s��"��IJ�N�Q9������وt����jVѭ@�y��j��kj�����N��L����͜�}Dq�f��5ߧE4��L�{	����Wma9h8wc������5���!�w(�y?�?�JY�)�Y`��jD4�7�癆cg���&Bzv��`f�(��H�RtV�^RD�+����N�ǁ�f�T��p_U
#��ʟ�1G@<�6�Q=ٌ�{m�tOIkV�g�ػF:7��*W�;֒	��x�(�6k�4d����Fi��I��RhF���9���x��
&\C��J_�0����O��Ě������������0u�\k|RSm�y��c!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc>sh�ڌ6�ve���'�=�9���bg2r0b�wa�!��@o����8����`4�+��+ER��{ia,���ߡ�c �ج�γI�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U���|K�{ߝ�Fc��B�I%ji�7��
#>:��� �rmd�&l�����i�I��M�3q��=$���A���ۖ?3�'����1Y�ΊS&nQ�rV�kV�џ�}$|~ïSup�xg쬉� }�A�%��fOX��8�r�;T3���/�"[Ʈ��JHn��z�F�x�aK�k��GZ>.�004@�k8���F�5/K �*jE|�ڴ�>��Xӌ��=)֞�)56s@��t�N�}�`�k��?Ŗ��R�A�%��fOX]a��1qh_�n�To�[�C��-��JHn��z�Lqܳ<��J*�Rs�0��(o <[J�	�LÆ�ѯ�x��yŮ���z��!z2}s�Uʚ7�ܩ�.fOe	Ln��S�W�"Lq�q/��Q��ǺΕE4���0Q��J���6�,A)�ؚ�����
��\�H��/Sg�w��'op�[�d�3���`�kq͠|�zDN�-�!I��'���N�"9���b�=����r{d��JHn��z��c�Bo��F:����Į��KH ��ߞD�ǒ�J���6�.X��;;"����v������*�%� �2S��(_�<��=k�Rm���Yci��zW�F:����Į��KH ����멋��I))����A�m�(��ʢ
w��]��0�ȍ�x�>c��w��'o�Q�kŕ��Q�Ӹ$P���F�׼K�3
�v�v-}�	mp̮�%I�����0i��Y��f������&J�b, ӫ/��m�B�K��1Ҹ�]��0�ȍ�x�>c��w��'o�<���q��q+����>(\�H��/Sg�w��'o�6���OB\�Ns&x������F�׼K�3
�v�v-}�	mpl�!����_�n�To�[�C��-��ɨ]^(���Ѹ���_�j�`���: ��ao.\C�k���uf|ò���
��_������B�K��1��n�da�ۣqM��X�~ ӫ/��m�D�K�h�x#�L_ѭ�Q�#3�d^�ϓ��ͬz�Ť��!4�%�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�oZ�o�S��	p���DUeH��lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL�t�� ���OgۈPML�����"{�B���}$|~Ð�BY
���wb�S��V��^��\i�ֱ�q������m�q�k�v_Q�(��Қp%�0�ΩyO^~�R���ce���n��8&���I���|I���:�Ϊ���L�8ɵ��i7N�_�M�3|r (���B����}�-�f ���:=��1���h�E)�.�2u�ɯ/wI���?����}�	76�&�R�Q���~��p���웂���a�"<b��5^,��*V�m��'��3�V2���i=�d����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�i/F@���V.F����R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
���y[6���ڀN�&jl�o2C�g�kgw�"��I��R� V�pFr����A"�U���w�c*����W"��ό���.�d=��¾ȼƸv��*Qxm�QA�Q* 5�����}Y�]��h@�YyZ��}�Q?M8�f2$ Hl�]��u3�0~͗��3��}�	76�&�R�V�"�0ɶ37y�����:��Y�g�f��߼
�dUY��~�6� ��5}�Y7s�9���o��S8��@糺뾃7܌:����3Eֱ�q������m�q�>1�Pq�@\w��0]���8-|�Dp��xs�S�)P<�ܓ�Y��=�g���>��8��-�Ϡ���:=
ҭ�3���VFc�B:�pO���w�_fHN��R��Gu�"�0�R�@�6�֐����o����(��e鎃9���1�L�]�b�֘m��+��$|��;D���J7"Sݠ�UM