��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�\�� ���K�O�{��?f���ʈj��U�sqc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<�w�>��S�Ś��
��H,7!!?�#�1�:�Ω��{:R;ޒ1 T�V	�tL��	ǖ|�NiUR!�`�(i3�q�9�ͭqt2�*�����-�/Q!�`�(i3!�`�(i3�1B��ӿ"#~j[O\�K�y؄@�!�`�(i3i��ԇl2�����Vc�r5�:�!\Vn�w;J��w�4
>2�����Vc2�����VcJ�g�Hغ!�`�(i3ؤ�$!Ѫ���]6'�u2�����Vc2�����VcS� ��y�t��|���2�����Vc!��.���j~����B��S3��V1֛s�ӱj���fI�i3�������8�e$�1�D���")�/K�L���\��2 ���J��&�S]���}��U��=�A�PvH���mwWA���c�0�9���K��S���9�Ec��H�>)67F��UH&��p�M��Z̸*�����&�SV��"����R�i�cC��D^W��|��0����WE��/���h��p�f"���r������4� _;��i�1],Aبs��0�}bک��?���)t��⫓���3B�Hj7�lu~�~�y�Ap�1�G�$U��Y��U�W�8=�V����8ɞ�mQ�Tr�>b�L]���}���h?���+�t���P�����-ӅC8J���_NUl��FC�쌓���ew2�\��M!�nz��m��+@ˏ^ow�Y�`�o`d�kN���9�ĒTC��0���M�<lbts�I�Λyi�ZN�x�w�>��SU��Pa���PPe7m��������n|s�)>E1&7W�$J�|(�����	x]�<��O~��������@���0f�*C�"�L��v��d���.���X�����]��#���X
� �AH�ah5J�M��
��m6g��A� �oQx?F#��_L\�Յ�B�֪��Gu���h}j����5T%p5U\�����	x]̅���OI�}c�J�M=�-ě��G�$�5�	�s+џ�_�v%�L��xE*?V����
� �AH���CdZ�G�u� �(��Z�N��\�T�ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P��\�4�s��u�@�
�ԟ�d[u����lf/����Sd,�ϱ�)ů*W.Ӻ�bl�k�]vX��J���{�Z�JQm�!=�y����h�}�)���32ę8�����8-���/���Sd,�ϱ�p�`����j���$5�?� �٠FN�[\�i�]|������)*�M�����V�^�&�����!ښ�m��<v���ٌʪY�����iUM?a9-�7-ڍ�qL�\�X���щ;�a�g&C�V8����0�P.!܃��L~΄gO�3�:M7bR�u��w)�S�5� �7��Mv�9*���f��^.Ğ�	џ�_�v%�>+�$�~G�6֜S��0 ��D�W��.~�٭�Jر�D�8�>+
� �AH�)��H�� �b5z��j1�&G��	�����ロ�*�T������|�OA�
܊��?Y2���3")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QLi/-�#���'p�@�I�?g�f���\X�<����8��U�w#���y�֑�/6K�RZ�NCIw4t�iZ]XF�������̇��� +��u*K6HT�����Np�S��<#l=���E����F�'n�^0o��~+�ݗ���3^�����n����\�v�e�g����\Y�4Eb��Y{�o��eŭR±���]SBÀcۄT�٥��T����kF����K�ca�?��J��Z\�'n�^0oM�D�;��-e>����C8�����M�g����!�`�(i3��|g�Y�'���Xw��������lԇ�-{�Y%T��BPe.��xu	�>��l%i�-ʲ��U�4�E����F��j���0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6����^���m���>!�`�(i3c��Et��q���U��>�w�Y�#� ����������5	���]���>����C��"��K��~f�[c��Et��q���U���
��I��N�Cٺ�������5	���]���>����C�/$�ߺ��]�P���Qi��(�
t�ژq���U�[��N�������l�
H�w���]���>����C�pॻ}��!�`�(i3c��Et�Y�{'%s��.|Z���ǚr��y�_��wBW��8���/�y����\mע������Y%T��BPe.��xu	�>��l%i�-�Wv�4�1�>��Z{����|g�Y�'���Xw�j�7��a(􆿳����^��/Z�o��>��Z{�Ǖ�(�
t��Y�{'%s�ui�铨g��U-�e�,���6+����3rn��yn_Fu��TD��ό���.�>�Q�c6�`S��|���Yl���#�]�!����M[��Ǣļ$����"�,�>E���TD��ό���.�>�Q�c6곍�ٜ�]Yl���#�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳����^��2�0���Q�#<4^���(�
t��Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9���6�e�:r�"J��M+7EEN�p!!v*!����a0��\�ټ�]�����q���:�0a�0��+3ǆ/������}	���w��Ot+�z��7G#+��\w��0]�m��
��1���&���]2�y�Z鎬���������o�	�*ZV)�J����67G#+�Ǘ0z�cUL|�]���?.�9$[{^7��y%%\�HP@�a�~�7���� ��JL�N{a�9Ow�Y��k��ı����V���}���s+���j�޺�5%q�P ڨ��S���Qߵs<��7�m��+�<4��ˌ�ň��h���T�%�/ң��Z����UV~s�"yp�m~|���Sf�l5/׊zo��'n�^0o�'vX[���am��	t?�*|�c���}i���o�dŚ1N�z ��y��G>u�\?���Y��i�s�����E�eNzL��<�7>!s���!5�e`��9nS�dB��,�:U�h���<��j����k��#�M/*�3���+��q2�C��i�j�kѶ���� �(�Mz�Iʬ�v�z��]'���Xw�j�7����'�\�n`��!��B�T�\ ��i3�|)sՀ�T�ya�����	?����n`5�fK�\w��0]b!��uፍo��ځס�^?���Z鎬�����}�f����a�Ň�b>�"B�ߋ�}�
�?�l\�=�]y�зq8�Ј'���Xw���,D}p$_~R��1�U���]�!����w�Հ�b02�O�.;}%;A�7s�9���o>��l%i�-5�e`��9Q�TyǨ�h�2�6�>*"v%)��2��������� +�ϖ���~v�@����gG���_����e޸XhZ'�kZ��w�rs�i�kۜ��/�X2�B���s�_��wBW��8���/����,D�C�:�S��>W�~������+�J���q���U��@����gG֫>����EN͞�!G�d�٣��c�A�L'Qī�*pY��am��	t?�*|�c��T�\ ��i3�|)sՀ��R�A0^L�ܲ�k?��i%Q,$'���Xw��9�"�5�-ďH�V��#��6�n`5�fK��0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6���2����.㓁bA��F9�0���ݼ}J�AZ鎬������_�,���t&�/s�2X��K����P;!).Y�{'%sAX���	q�KS���K����)��T�\ ��i3�|)sՀ^X��:��h�b��0���������q���U�h}Nw���M��_e޸XhZ��Q]� _�rs�i�kۜ��/�X2�B���s�_��wBW��8���/����,D�����ߨ�����`�d�٣��c�A�L'Qī�*pY��am��	t?�*|�c��T�\ ��i3�|)sՀ!���fxoo�c�S��bƲ��+�J���q���U�Z��O��<�"��~Ǣ�)�s�ި�b!��u�[��l�,n*�"gg'���Xw���,D0��R�iF�h4M&Y<1�d�٣��v_���Zo��u��Y'G�7s5kL��d�٣��v_���Zo��>D��e2���HF3}�
�?��&��>�!�`�(i3�d�٣���N N�S��30���,"�x|ٲ�зq8�Ј'���Xw���,DH�v����ܕz&�8�n`5�fK��0z�cUL���.�1�3�8���/����,D�x ��s��q���nm�n`5�fK�\w��0]b!��u�s�Uo���]H/��d��]�!����w�Հ��}�a��>�A�IS��#�$�~�M�q���U��@����gG5m�E��P����z�7s�9���o>��l%i�-ݓ��E�1�#��d_�E����F�'n�^0o**�ХM
�nGZ��JP�O�?~Gv �@����gG�S���!�`�(i3�b9����U_�+X�Ă�L�i�;#�����v��#;�7���c�t}���#���Q]� _ό���.�}�
�?����S&�r=�������d�٣���N N�S�+w�7�
�p�	%6зq8�Ј'���Xw������LƑ���@�&_E�EYZ/�+V��i|���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�"��B9�
eBZ�tX ��Dsa�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WD�K[�,�ᖠZ�q�PO4�7��V���.g"}�p��q����`U��:
1������Q>ml��B<�D-��I����~u���3rn~{�3�����w���H��(6��W� ��iE��lN���2�0����(@CPw�>1J���Va�%��jqm�
���n�ѩ)e�qjn���H����/�;�ƽ�/��e޸XhZ��_�#�:�b��tT�ę_A�7�UyR�jt�Q�S�O�ώ[���ػ);��AY*�Ld�!�`�(i30����3�0����%�/ҁ��:J�a$�Y ��!=w�- �n}沁2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �O�t�&~f3��gL��_a;�+k#QXO�S�p��QM��b�(�2ɒ�E�-��%�Y8)=���a�Ň�b���Z����I�>�>�F�1I!6�xˮ�U3޹�:^�a�%-�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �*�<��"�U��)���Y;e�iKI/B޾Pb�i0[����8|bs��2[�a��o���H�RtV�^�Y���GiL�~�*qA����6\�4�@�� �-j�1tSjv������_�l)����Aɠ�T�nGHN��R���ء�I��߸��S�Ȍ�b�W<_|���s���>��FS&'ב%��iK�D�b=.��6��=�Y��q�$���t�T�ZL���hs��>1J�����1�谏8Ҫء�6QIl����!�`�(i3!�`�(i3��A��
r��G�
�M���)Y��"����Y;�"�ff���Q����(�u���ݚ�Н�!�`�(i37�wtMMJE\&
��d�G}%����3f^�#Ҧ��>-�`<�K���$�N}ܐ�E��D�G�&ց�*�0$߀���9��n�7�Y���_j�����9�x�\M�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^�Jo���jk���%�8�Va�ir{��b�b�*#o�]�ʄ�v�4�?zm�jd7}�� ��M�sv��>���F*G�D����ݚ�Н�jCH�d*��=����h��LAи�!�`�(i3�I��Yqt��ۻz�˾ �����]M?��y�!�`�(i3m�����G�FW�DVx>74/���j94�JW��
�:qEp'{w#/ B!�`�(i3��w�`L���ǚ����}Dq�f�HN��R��bP�63Z�t�߆�p�h� ��5%q���f�e�&�U��f�!�`�(i3�FW�DVx>74/����j�����HN��R��F F�E̠(*�O�q���}���wCH$�I��*�M/*�3��q�t	<!�`�(i3����,����0�|�_�mS8<�n�ݚ�Н�X19�-.|}�ڎC�?�x��w����/�dI{�b~*��s��J�'Ƕ.(�����1�OG����ֺq٫[_�mS8<�n�ݚ�Н�jCH�d*��=����h��LAи�!�`�(i3�d������7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j������
C�ݚ�Н��̢k��� :b/�Ti���i��1tSjv�!�`�(i3����-Jg8�iT��*�����B�fĉ>99��A0ok�Ra])n#����,����0�|��';��#j�ݚ�Н�-��)'�>���F*8k��.ͥ�H�RtV�^CH$�I��*�M/*�3��7ݽ��!�`�(i3�k��^�1lv0�9l�'����u��r��!�`�(i3��w�`L�P�~�9��}Dq�f�HN��R��bP�63Z�tHN��R��F F�E̠(*�O�q]q�iE�>�CH$�I��*�M/*�3�F�N��9R!�`�(i3����,����0�|�_�mS8<�n�ݚ�Н�X19�-.|}�ڎC�?�x��w����/�dI{�b~*��s��J�'Ƕ.(�����1�OG����ֺq٫[_�mS8<�n�ݚ�Н�jCH�d*��=����h��LAи�!�`�(i3�d������7s5kL�G��Hb� h�ҩΪ���l��`4��C�<�5��t�1tSjv�!�`�(i3O8��u��8�=����h���7�)��~!�`�(i3jCH�d*��=����h��LAи�!�`�(i3��w�w:�!�`�(i3CH$�I��*�M/*�3��q�t	<!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN՝� s�#�=�U�u�íN=]8k��.ͥ�H�RtV�^pT/�GS�7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j�����>�nE�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub����pT����d#��N�Q4DҚjjCH�d*��=����h���7�)��~����l�� ��5%q���f�e�M?��y�!�`�(i3�%�r����ֺq٫[_�mS8<�n�ݚ�Н�jCH�d*��=����h���ʘ׋�\!�`�(i3�I��Yq���k$ ���y��lD:G��}�/��f�\%��1���g!�`�(i3���F��O��ݚ�Н�T+���f�ԬQ���Kͽ<\��1tSjv�����l��Cd��9s��vr5�Dѯ���-����!�`�(i3�FW�DVx>74/����j����ʉ��%>�rGO�D mWN���%>�rGO�D mWN�mJ�0�6�ʁ���Mյm�����!�`�(i3��w�`L��^��&vb��}Dq�f�yhޖ�k�j:��e+�������� h�ҩ��H�������+1�;�.��1���-����!�`�(i3�%�r����ֺq٫[_�mS8<�n�ݚ�Н�9��n�7�Y���_j�����9�x�\M�ݚ�Н��Ra])n#Y�5�n����N6�������&G!�`�(i3�� л��OP�Յ��C!��AVt���r����Վ~RT�ط���RƝ"�f1e��&� ~P
W!�����T���ݚ�Н����y��lD�ԄQ/	D��p�����E&R�v����f���1=ƌ�F��ſ�c�<�y�u��!�`�(i3�FW�DVx>74/���S�%�[!�`�(i3�5ߧE4��!�`�(i3�k��^�1���+1��*Hx�g���-����!�`�(i3_��5��p���E{�ς=I����`��"!�`�(i3VZ�ڋ���Y���w2dv)�
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W���	�N�M��/�9ސtjCH�d*��=����h�TGaG��7ŕ��aR�HN��R���
�Ŏ����ܐ�}�^�#Ҧ��Uw:����/$�ߺ��]��6�
V���M�{�|L�8�YX�s�m��P4-BKI�^$D����[�#�������#��[��o}�	?~h���X��*H<%���!j������,0Y�z���h�
nЯ�O�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3ޙp����ԬQ����5��t��}	Vӯ)�^C���r�/��tM��� !�`�(i3!�`�(i3�>d�g�K���S&�r���d�L���!���乍���Tj'{w#/ B!�`�(i3}Y;�jn�Q�rV�FZ�_v(��ڥ����ȾrB�WD�{����0��e���F�&����N�='{w#/ B!�`�(i3}Y;�jn����>�~:w��="P 2`�����t�ؚA��p�W���=+XR _;��i�1QR ƫ8��K��6��@���ɗ;�6�[�:W�N����%{�O<���1ə�*!��F)_8���S+0sYҔs�8��C5W��W�݈��0����=sv9jV Al��4���Ҧ��f�F��(�[�o��_�Rv�䩲$���dS@Ɵ�o��èVxjzӝ���I(͂��-����;�~��-�f����Ga��'DV���b�z'hۉ)��d�7�qĮ̢k���F�KD�Vr[/}>5��0�B� �b���H����@��	Ķ=��h��t1p��5�F���0�|�9�]��۠7s5kL�eW���Z���
nЯ�O�f�"*&�k㎺�s �Ա`E�p����S{#�lܵ�"ǉ�t������z���B� �b�Ъ���l��(�Mz�I�-Ki�\�I� �����;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���wFB�b���\��-&�C�U��)���Y;e�iKI/B޾Pb�i0[����8|bs��2[�a��o���H�RtV�^%w�*�7��E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��c5ew��ԬQ����5��t�	���QC�꠼*d�m<���H1tSjv��H�����3i��U��a=j��� !�`�(i3h�@�F��:�8QG8�]߸��S�Ȍ:�^ao�a%��w�ݚ�Н��V�qZ%	L:�U��!��(�Mz�I�y:�1^0lf՝� s�#���k$ ���������'|Fpॻ}����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�ȌM�����UT�GP� �&���N4����j��T6�o8:4�I���c�90��G��6�iI9�o«IX0F�M���3rn���Z�[�[�'ž1�|�'����u��r���}��C˥�!��_�*9 ��b+}y[�k��^�1��dc�@c�����h��-����J$�,pW�ԬQ����5��t�;��Cٯu�Xy|�W1F#�֞q|�|�������t��Һ'��b���͵H�L���j#o�]�ʄ��.�L��w)��
=b~*��s�l\�=�]y���4y��ij��X� 2ޙp�����,�,&��`�2,�!������������xQ��
nЯ�O�A/��M����,�,&�u?N� ;0a��>L��,:&Ȍ�g�F��6�o�B�Q�BB��A�^f��[�#��^����B.l\�=�]y�z���^F �K�Ǔ�\� h�ҩζ[�	���d�~{��#o�]�ʄ� �
*|'pUÉ�L�XG5���Z/�&��o��4P����9-����yΪF!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�U��ýPe�O��Ϡ����Yk��1���~m�ڨ�hծ�d�tuѩT��Z|�����{���}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�I֬W.�dD�%���o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ܝ�s2���lI�k4.��7�t�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�TM�a��G��P����U��)���Y;e�iK!���d.���+�^n=\f�5>���௧��T×r���"sS<�0�zG�������&G��������O=�W��E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv����q�D�-c[����dN�<@Iv��nt=:��:5A��p���KL���>Ht�u�UG��Hb� h�ҩ����q�D�-c[����ӲY����&
@!˥�I:��q��k��^�1s�Uo���03�� <I�����&G�����$ZtgQ�9OZ�s:�8���Ӫ�Ġ�9�C�s�4՝� s�#�,��&5d�:�.�N�Ĺ�Z<��A!��-�����d�tuѽ3y��;��"?��FZ� d�!y�b�G2fĉ>99��j���Gp��Ě���aT��3G�IX0F�M�27���^��~"�KT��+Y�6R��M�,!hޖ�A$�P������5d��n4s1�U��B��-��8�2W6��v�����r$ɓǃl[�Ƶ�1tSjv�� �@[�鋽C�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩξK�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�irD3w��'��a��o���H�RtV�^$����}��*�f;��}Dq�f��5ߧE4��;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���r5�I��drB�WD�{����0��e���F�&�?\MP!� u��r��J>zߋ��>ַ�����ƍ2���l���Ě����E�i�m}6O�D mWN��ܐ�}���$�uG�N6-	��6<���oA�LD!�GkǤ661��������C7@�����hH��6�3��N�߿�wW��ZN����6�o8:4�I���c�90��G��6�iI9�o«IX0F�Ms�Uo���ci���{2�'ž1�|�'����u��r�吆v��7�tG��!̒j���b+}y[�k��^�1��dc�@c�����h��-������Ϟ4�>Ht�u�U%��v��;�jmT�#�0M�Ŷ�Eʨ�`N/�a�	�Z����ڎC�?�& @=F�S���iﳣ�N���V�Ո���߿�wW������4Yz����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�m`����Z��b���Q>�<��#b�8��B�5�¹�*��a"N����#�T������oj������ZN����6�o8:4�I���c�90��G��6�iI9�o«IX0F�Ms�Uo����=Djw�9�xjzӝ���I(͂��-������Ϟ4
T�W��%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<Dw\����ō܈��VW �+��}Dq�f�����,����0�|섃Va�irƦo�
�ƳI�^$D���5i�a�vb�(���27:�������&2��OY�J�M����!�`�(i3s�Uo���[;\v�a���?D�8����Ě����E�i�m}6O�D mWN��ܐ�}ĚȜ��Y���܆��줬;}it���U�R'�˴$�#��Q1�dfC0o�4��F�悠A�,��b
�C�&`�@|�v��������U�Rdd@��2�M�,!hޖ�A$�P������5d��n4s1�U��B��-
r�	O)�A�IS���=Djw�9�xjzӝ���I(͂��-����w-)Sz�M�:�.�N�ĽC�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ���U�R^p���P#%��v��;�jmT�#�0M�Ŷ�Eʨ�`N/�a�	�Z���Lm�<o��!\��� fa�н(�P"G�wk���zܳX�P��%�©��-/a8X�o|3bK�����`���UK�"��ӌ�rHN��R��bP�63Z�t�5ߧE4��Fr��jlk�p�+N᢯��0��ĥ�A�)�'� o�F��(�[�o��_�Rv�䩲$��8��I�:Fa�7��׏�������u��0C�r$ɓǃl[�Ƶ�1tSjv�ٮOS���p�]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����-����;�jmT�#*��m�vэ%�K��^/p#��I2�8��[�@��W��*����!�`�(i3,��B�u���Ӹ?]qt���-����!�`�(i3��S�V� h�\��;�,�Ra])n#���r������!���Ĺ�J�E]�?-O딈pᜯ}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��{+�t��Rz�R�k��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�sݸ�/�gxjzӝ���I(͂��-�����d�D��^օ?D^���k��^�1��dc�@c�����h��-����pT/�GS�~�+yp�l�����z����-����;�jmT�#<��4�e�AԢ�a\�2}$#h6��8{4����g�B� �b��!�`�(i3�j<��?����"���w�w:�!�`�(i3u�st�⫴�IV�*F/��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��̓-���.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc63ͼ�a+��X�\�[2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�"�_�Ȫ��q;�4���W�&]�6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&GZ��JP��V��#��6x����E2b�z'hۉ)��d�7�q�e�OB]�4<W��Q��ic)�̩ƍ2���l�;Tti�����|�g�'DV���b�z'hۉ)��d�7�qĝÜ�f��E�h�b��0S^Գ3���ƍ2���l�����g�Z��3��a���!@�f")u��r���\!�U,ܓh�,��R��3��
�M����d��-��!�"ǉ�t������z����-����H������N����ӄhD����6�i�|?���S�!��EF9�0����ۏ�:��"�vW(�����C�Y�\�=�40]���8�C�Ћu���ܭ i��h�
d���@��3{5�,#&WJ�z�6�2�^�?�.g"UƄ3[�g�DPp���Ě����E�i�m}6�@�	���Ĕ׹�4��)'���y�Pc�1�5;�����>2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc68�=��l�`s`�� �n�җ52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�D��Ø
���R>��6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r���D��Ø
����vۂ�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK���7�^t��d��-��!g��J�s����0�|섃Va�ir[��l�,t���H[W?G�\̒=��3��0��{��b�b�*�,k!��L���Vy�`��vN�[���}��W��L
��r͞�%� h�ҩ��m��
��:�'�:5�y�����;b�-�2��z*	��y��R�o�"c�Pd�BR�~;�A*8k��.ͥ�H�RtV�^�D��Ø
����vۂ���QЪ��\O`�� \)���F��O�}�	76�&�� Ӗ�t$�)�vx�ӽg_ʇ4�C[�#2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��z��w��N 	���;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �n���H�g������φ��<�6�@a� ��fFMqlg��èVxjzӝ���I(͂��-�����9lD��XH�ܲ�k?�#QSU:��8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�D'm�����Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s��ݚ�Н����V[���*φ�\-�gM�?L}�7�n��<f��5p�T����՗fc<1tSjv�K��ft����Y�b���v�Ѭ������:t����0`T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH�ܲ�k?J.���\f��V|Cq��Ɨs$f��_Ub��7��G_���;�P�t�5�׹�y���3wϮ�Y�b�κ/^a�_2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�{�ը7tW�o&w&v"3��?�32�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܺ�5�������@����	�Qߙ���O;�
�,I�@�"|�n|s�)>o�oNS�'Y��s�_}}
�;?�c�@��B`���~��~\C�~��/�T�٥��T�5�Y�w�� ƈ��V���TtU��
�IȤ7�����t�T�-g�
M��Ն��5(&�L�����Y�z0=�_���{_8�Y��=�}�Vݨ��Qu���%y����c�S�ڬ��M� ����%��ӟ�u�g�ly���
��Q?M8�f2]�Q�&��H'o�a8��v��ONH!�`�(i3i}B2>�~ �<j�"�AM?��y�!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H��Ⱥ�Q���'g`$�YD ��� ��?D�8��HN��R��bP�63Z�t���������l��Ht5�=�5����������&G!�`�(i3
/���p\"�!˥���KS����<;�$��\|����=�'�^�����ݚ�Н����F��O��;b�-�2��;�P�t�5���W0�]ݽJ/��v�$�)�vx��ef?���Y=	<��Ғ*H��M�$��ꤹ"�ۨ�%�ۥm�Z�]�.nŕ��v��i���Cb�Lc�^[v�58u��\quA0�e]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^<���d1x��r-�TE�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t�	���QC�꠼*d�m�d��-��!|�|�����@��pr��4N�J�ף�<Jq�Z9��5p�T��e����[�v�4�?zm�L�[\�"�B� �b�ПB�'��a��*ZV)�J3'T��߷j��
��e޸XhZ��}Dq�f�m��;���1&��*�("��X2��4�j:��e+�������� h�ҩ��m��
��0: ��q��%��j��e޸XhZb	�fƏ���%>�rGO�D mWN`���*1���F��O�\E�W��4b����A��c�^[v�58u��\B��U<2+#2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�*I��A�*u�>cC=V�g`P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc`��P���P�L29:(�U�E�0�IDKO��	h�{��-�wXB`d����3�#quA0�e�&=u������FmvU����èVʲ��U�4�a޵��	dN�<@Iv��nt=:���2]���`,9�H�W�0��K�[̞��>����� +"�*aPV�6�����Q�8�w�[���:=r��Ɉ�?����2���-/a8����l��Ht5�=�5����������&G!�`�(i3��	~r��k�%�D����MxOܳ����|e"��w�w:�!�`�(i3ʲ��U�4f�
"_��P��]�/F�ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6�E`����Fr��jϤ�LǀN���)��%A���h����u|�
�xr�{���г��r ��T���yo��5�I�B4�٫IX0F�MV�ҁGG%4vkz����`���φ��<�6���w���c�ShT���A(�c���_G��Hb� h�ҩ��W� ��iE��h�{:m��b+}y[�k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vNd�8��k�Ss��Zf���g�F��6�	�¥�S`Q�TyǨ��&��I��"ǉ�t������z��rx�pj�d�B�'��a����w�蓺���pJ5�!����;b�-�2��z*	��y��R�o�"c�Pd�BR�~;�A*8k��.ͥ�H�RtV�^�<��a�X�r��ڵ�r��@eM�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b�[�؟�-��@뀗2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������y�$��_,�����{S�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc7=�� C7<;< }>�5��Z)l�<#l=��,�W�8"M�5�O�%E#PMQ���0�+ʛ�����'�PD�{��b�b�*��ic)�̩ƍ2���l�=7�7K�P�"ª���aT��3G?�d���&��]y�Q�';��m-�/v7|�|��5��Z)l�<#l=��mWᅫw��K���'h�x��JyKc>�9k����ǃ_7^�	������+˃��ƚ��o!��yV�oD���w	����hz��w��ￓ�����J�'Ƕ.-�DAԄ��'�i�*ڶ�UKs,��#��I2�8��%��I���L���͛|�u�ݪG�B�	z�W��7�3Z��ȍ�c0B�:
��t(p���}ƿd���O�&s�6q��f�,�k]���d�L�ѱ���F��k���%�8�Va�ir���+1�;�.��1���X2��4�j:��e+�#o�]�ʄ��O��:���� �!�ա{�4����0��e���F�&���J�������u�h1����jd�	�!�`�(i3{�d"���毘3)�:�4�5�$��GW���6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3=7�7K�P�"ª�����}Dq�f�����g�Z��3��a���!@�f")u��r��;�E����0|�mll6pe"}��\*�>1J���KT!��ĭ%���G��_��	���}�J��"�W� q��j�J^�G��
Z�g^!oA�Pl:�����Ǐ˨�g����m�5h1���'���C&b~*��s�φ��<�6��`䘸�|������&G!�`�(i3	�%��6� ����7����|e"�̢k����m���>#o�]�ʄ�M��,����q���f�e�G�\̒=��!�`�(i3�{3��������� �!�ա{�4����0��e���F�&���J�������u�h1�"�Yt�㝌b�Bϱ��e�P����E.��.KV�9\�hF
FB���ՇdH�RtV�^�i+��9�̪=���"��ӌ�r���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�~(������
���F�<��}�u�?�d���&��4�5�$YA@�H������f�6���t�T��?E-h��`f���sd�G}%����3fJX �����P�2Hxjzӝ���I(͂��-�����i+���c�1���7ƍ2���l�����g�Z��3��a���!@�f")u��r���m�5h1���g�F��6x��w�����ԬQ����5��t�	���QC�꠼*d�m�'����u��r��i+���c�1���7�?D�8����Ě�����}Dq�f�N�-�}q�0/0`9N1��-�����#�-�p�%��a�����b+}y[HN��R��bP�63Z�t�5ߧE4��Fr��j�p���"sH�",r'�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcU5.���}���\-��U��)���Y;e�iK!���d.���+�^n=\f�5>�.F<!W��ShT���A(�c���_G��Hb� h�ҩ΋�Q7lY��״$(�>g��̢k���F�KD�Vr[/}>5��0�B� �b���H�������3rnu�j�fK������&G��+�t2�������/��kOT$f��_Ub��7��G_���;�P�t�5�׹�_S���\���{,�M�|�Z��T���e����H���,>$��:?���