��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��]	h8��`��(	�t� �c�=0N���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:�k��X�.��ѫ�� �mD�?ea�8���`8��xS��������]P*m����)O��Ξ4�"�\�� ���K�O�{��?f���ʈj��U�sqc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c,� � U�rN�3��m-�@xI+r�� 0�D�A�f�mX��VNF��SK��1��sʕ��͛E�{�ڌ�2���2��ds£����&��ea�8���`8��xS��������]P*mQg�@zh�S҆�|n����Շ_ Q �y�N��Q(�V͆J�Й�m��x����y7���̖�}�Ϫ�h�C �@nk����k�&�J���qݣ��6Q�eѢ��x��!�v�j�|�㈱�U^��\�4�s��{��]Qǯ������W)����VIW	I��?G�~�MUs +������\���T��U	�1�_u���*����	�����	����LO9� �Ŭ��2Dm�x]��.] �'9�����L.��6�H�.���2/�f��=V"N�^{")8�*I�ց��6 �����Y<�zd諒~����L.��6+Q)?^R7D�y�B.h�hC���(:�J�5`xt��R�/E�CԵ�_�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_��c�W_QL��[�nh�/;KYˆz}()pxt4���J4xʆ)�-E����}�����b���q���1�:�Ω�S�T�;Ϗk[�^��_��c�W_QL��h]��������@J
A��w|�<��'p�@�I�?g�f��u�H(�3$������/�����,��B	hI�ˋ���p�ϵ�DE�U���JHn��z���G7���}9s�X���@�X��l0��F��j�q	k���Aj޽���Ǜ������`�����"IÙ=�H<z,Ҽ&�כ��pܔ��n����\�vņ�Q�]����O���R�^Ƒ��l0��F��j�q	k���A)٠���ٴ�]c���HQ�n���{�)w�<�_NOnRI���meo����\G�Y����-�,��Lt�2�t"�,�>E����-��%Mό���.��_F�k-�!�`�(i3�����5	���]���>����Cοƿ�d���!�`�(i3��|g�Y�'���Xw�4��}�<������Ə+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�Hᴕ��U��5�%]���a(􆿳����^��u��g��L�������|g�Y�'���Xw s4S�'�i��`�z��GZ>.�0wa.X�wY�����ϲ�CyW�f�tR�wX��q�\E��0	ozqP�"B��$I��w��,�������ݹ�0�����иܖ��+V.���W����vcy��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+o�Tku�����F�N~Y��C�Y�)��NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��u�H(�3$������/����5���N�.�����	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�B'�P���i�(�S���N�؆�B��W+`�x�oP��@t�&�e�5
��Ib����rs�i��@�N3,(�����ϲ�CyW�f�tR�wX�����/��&/9[�L\����	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8��H��rR�^Ƒ����"X��[��Q[R�7����$�1�������7��Tl���W+`�x�oP��@t�&�e�5
�\l�'$9��`�[�*!-R�^Ƒ����"X��[�d�a�4$�b!��u��<��>���%�-�]�Ǣ�V0d%{�;����f�kN�ı&l����[}�@��L}�
�?��u��g��L(���x͢'����&���Z02��`�z��GZ>.�0�i�ܰAb!��u�\.�l������^�i���"<璋���n�4�{lGD�V�B��иܖ��A�.u�rI����"��T:���V������?��O�/5�؀Ǣ�V0d%{�;����f�kN�ı&l����[}�@��L}�
�?��u��g��L���NE!/�3$�+?>5ܔp�l
d�R�.��On��M��ҹf�f3'i3�|)sՀ�/V����!�`�(i3���^��������KqZ"�V�踫g(�r� k�|6�8�S}�3�U����.���nH9�ئR'cf���a�	& ��?�d���&����]�p��>�n��-ؐ�	}�@�r�<Uee�,�Aٺ�H���H�V�����ѥ�)C�G����]'\gWg��	�Z�kfc��2���8���8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�?KYC'v���ʗ�%����صW�my$�N��o�/���;�B�'��a� 7�J�[|�m�ߕ�E�g�������(ӈ���m�r����m�ڨ�hծ�߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3?KYC'v���ʗ�%���S�*(�����Ə!�w(�y?�B�'��a� 7�J�[|�m�ߕ���DKY�������4�:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6���%5)R����,�ǰ��i��W�o_aP6r�ut�0o��F�5(��~�q��a��Se�������,�_--���g���R�?KYC'v�����p�*�u��g��L���NE!/������D�i=�d�w�R���y���,!���wMn����A�rD����}��\CB��u�Y�KG�	�v�3� k�|6�8��:�EB�Z5�O�%E#P�� ��φ��<�6�@a� ���N���������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�-��ټs�  ����'K7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���Pi�#��R;�jmT�#ފ�����x�Bi�v�V��	��7^3ZiY!�`�(i3�/�cLbŪ�����:Y�{'%s��v�9˞�]v1�_ُ�����Ə?X���V4&�]Pn��J�:�_q�pWS�*;q�=�9��tsȸ�"rR��w�w:����Fz�8��;Yv^�-w2M#-5�]�!��	Ǹ�y85��X��I�ՠ��t����>3���w�@V-���,W��AԢ�a\��MԵ�x3���ʗ�%oc�����!�`�(i3��Ě�����}Dq�f�FwZNE�&tS�D�]v1�_ُ�����Ə?X���V4&�]Pn��J�:�_q�pWS�*;q�&l�p�q,!���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}���L^-a�aT��3G?�d���&� ��G����8�C�f�F�5(��j���rz+��bc�n&��<v�\�b͐�	}�@�r�<Uee�,�Aٺ�H���H�V�7�}�!��q�(?��q���t�T��?E-h��$^(?��"��K�����8-|�D����l��A(�c���_G��Hb� h�ҩ�?V��j�c���o���T�{_8�Y��=�}�Vݨ��}Dq�f��k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��H�����Yu�������&G!�`�(i3{k�h�+&tS�D�'���Xw�j�7����rF��8ל�}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Fr��j��;������/X� ��I��)���W�w��fDl�s�K�6j�"Hs�X�8�x T_&"��ߦ�A���`����oȺf��m<�E��?�d���&��8� t>K]�S�^t�`,9�H�W��<��Y�&l������8y�Ɋ����Z���2��}��1�O����!���c�A�L'��b���A�&vY��;�w�R���y��E ��M�]$>A���w�R���yWp�K#J��_v��0!�FX���v�\�b�U4��\w��˪?�-���ei�^�̷ؠJ��:����}V�)c�`j�Txk^��]��3R��������Vo[���˚����Z���2��}�������Ə�m1�ؓ� ,��rQ3���w�@VeX�P�+$r�t�}iV��	��y�� �P�qN#?
]w<�h��R��e�j�Txk^�a���~6�z�����ϲ��Vo[���˚����Z�ם�.J7h��r��H�v@W��}�������D3���w�@V��B|_��j$r�t�}iV��	��y�� �P�qNy�WE~�YV��	��y�2B��$X|,�E_�CR��L(q_҂T�q�w��/��=��K�E��{#6�a?�d���&��D�U�2Y�Xe ��g[���K�J��]��m�;�¬pX��D�P�E6�k��q��־�W+��W�2W���R0_.��45��LҺ_.E��p���V�$r�t�}iV��	��y�� �P�qN�/9ݦ�����,�ǰ� Ϳ�&�vDv�}˨�� a���#