//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2012 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_SS_OCT_SOPC_burst_0_upstream_module (
                                                                 // inputs:
                                                                  clear_fifo,
                                                                  clk,
                                                                  data_in,
                                                                  read,
                                                                  reset_n,
                                                                  sync_reset,
                                                                  write,

                                                                 // outputs:
                                                                  data_out,
                                                                  empty,
                                                                  fifo_contains_ones_n,
                                                                  full
                                                               )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  3: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  3: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  3: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  3: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  3: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  3: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  3: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  3: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  3: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  3: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  3: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  3: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  3: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  3: 0] p31_stage_31;
  wire             p32_full_32;
  wire    [  3: 0] p32_stage_32;
  wire             p33_full_33;
  wire    [  3: 0] p33_stage_33;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_18;
  reg     [  3: 0] stage_19;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_20;
  reg     [  3: 0] stage_21;
  reg     [  3: 0] stage_22;
  reg     [  3: 0] stage_23;
  reg     [  3: 0] stage_24;
  reg     [  3: 0] stage_25;
  reg     [  3: 0] stage_26;
  reg     [  3: 0] stage_27;
  reg     [  3: 0] stage_28;
  reg     [  3: 0] stage_29;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_30;
  reg     [  3: 0] stage_31;
  reg     [  3: 0] stage_32;
  reg     [  3: 0] stage_33;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_clock_crossing_master_ddr2_m1_to_SS_OCT_SOPC_burst_0_upstream_module (
                                                                                           // inputs:
                                                                                            clear_fifo,
                                                                                            clk,
                                                                                            data_in,
                                                                                            read,
                                                                                            reset_n,
                                                                                            sync_reset,
                                                                                            write,

                                                                                           // outputs:
                                                                                            data_out,
                                                                                            empty,
                                                                                            fifo_contains_ones_n,
                                                                                            full
                                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_burst_0_upstream_arbitrator (
                                                 // inputs:
                                                  SS_OCT_SOPC_burst_0_upstream_readdata,
                                                  SS_OCT_SOPC_burst_0_upstream_readdatavalid,
                                                  SS_OCT_SOPC_burst_0_upstream_waitrequest,
                                                  clk,
                                                  clock_crossing_master_ddr2_m1_address_to_slave,
                                                  clock_crossing_master_ddr2_m1_burstcount,
                                                  clock_crossing_master_ddr2_m1_byteenable,
                                                  clock_crossing_master_ddr2_m1_latency_counter,
                                                  clock_crossing_master_ddr2_m1_read,
                                                  clock_crossing_master_ddr2_m1_write,
                                                  clock_crossing_master_ddr2_m1_writedata,
                                                  reset_n,

                                                 // outputs:
                                                  SS_OCT_SOPC_burst_0_upstream_address,
                                                  SS_OCT_SOPC_burst_0_upstream_burstcount,
                                                  SS_OCT_SOPC_burst_0_upstream_byteaddress,
                                                  SS_OCT_SOPC_burst_0_upstream_byteenable,
                                                  SS_OCT_SOPC_burst_0_upstream_debugaccess,
                                                  SS_OCT_SOPC_burst_0_upstream_read,
                                                  SS_OCT_SOPC_burst_0_upstream_readdata_from_sa,
                                                  SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa,
                                                  SS_OCT_SOPC_burst_0_upstream_write,
                                                  SS_OCT_SOPC_burst_0_upstream_writedata,
                                                  clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream,
                                                  clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream,
                                                  clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream,
                                                  clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register,
                                                  clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream,
                                                  d1_SS_OCT_SOPC_burst_0_upstream_end_xfer
                                               )
;

  output  [ 29: 0] SS_OCT_SOPC_burst_0_upstream_address;
  output  [  3: 0] SS_OCT_SOPC_burst_0_upstream_burstcount;
  output  [ 34: 0] SS_OCT_SOPC_burst_0_upstream_byteaddress;
  output  [ 31: 0] SS_OCT_SOPC_burst_0_upstream_byteenable;
  output           SS_OCT_SOPC_burst_0_upstream_debugaccess;
  output           SS_OCT_SOPC_burst_0_upstream_read;
  output  [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata_from_sa;
  output           SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;
  output           SS_OCT_SOPC_burst_0_upstream_write;
  output  [255: 0] SS_OCT_SOPC_burst_0_upstream_writedata;
  output           clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream;
  output           clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream;
  output           clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream;
  output           clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register;
  output           clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream;
  output           d1_SS_OCT_SOPC_burst_0_upstream_end_xfer;
  input   [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata;
  input            SS_OCT_SOPC_burst_0_upstream_readdatavalid;
  input            SS_OCT_SOPC_burst_0_upstream_waitrequest;
  input            clk;
  input   [ 29: 0] clock_crossing_master_ddr2_m1_address_to_slave;
  input   [  3: 0] clock_crossing_master_ddr2_m1_burstcount;
  input   [ 31: 0] clock_crossing_master_ddr2_m1_byteenable;
  input            clock_crossing_master_ddr2_m1_latency_counter;
  input            clock_crossing_master_ddr2_m1_read;
  input            clock_crossing_master_ddr2_m1_write;
  input   [255: 0] clock_crossing_master_ddr2_m1_writedata;
  input            reset_n;

  wire    [ 29: 0] SS_OCT_SOPC_burst_0_upstream_address;
  wire             SS_OCT_SOPC_burst_0_upstream_allgrants;
  wire             SS_OCT_SOPC_burst_0_upstream_allow_new_arb_cycle;
  wire             SS_OCT_SOPC_burst_0_upstream_any_bursting_master_saved_grant;
  wire             SS_OCT_SOPC_burst_0_upstream_any_continuerequest;
  wire             SS_OCT_SOPC_burst_0_upstream_arb_counter_enable;
  reg     [  3: 0] SS_OCT_SOPC_burst_0_upstream_arb_share_counter;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_arb_share_set_values;
  reg     [  2: 0] SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter;
  wire             SS_OCT_SOPC_burst_0_upstream_beginbursttransfer_internal;
  wire             SS_OCT_SOPC_burst_0_upstream_begins_xfer;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_burstcount;
  wire             SS_OCT_SOPC_burst_0_upstream_burstcount_fifo_empty;
  wire    [ 34: 0] SS_OCT_SOPC_burst_0_upstream_byteaddress;
  wire    [ 31: 0] SS_OCT_SOPC_burst_0_upstream_byteenable;
  reg     [  3: 0] SS_OCT_SOPC_burst_0_upstream_current_burst;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_current_burst_minus_one;
  wire             SS_OCT_SOPC_burst_0_upstream_debugaccess;
  wire             SS_OCT_SOPC_burst_0_upstream_end_xfer;
  wire             SS_OCT_SOPC_burst_0_upstream_firsttransfer;
  wire             SS_OCT_SOPC_burst_0_upstream_grant_vector;
  wire             SS_OCT_SOPC_burst_0_upstream_in_a_read_cycle;
  wire             SS_OCT_SOPC_burst_0_upstream_in_a_write_cycle;
  reg              SS_OCT_SOPC_burst_0_upstream_load_fifo;
  wire             SS_OCT_SOPC_burst_0_upstream_master_qreq_vector;
  wire             SS_OCT_SOPC_burst_0_upstream_move_on_to_next_transaction;
  wire    [  2: 0] SS_OCT_SOPC_burst_0_upstream_next_bbt_burstcount;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_next_burst_count;
  wire             SS_OCT_SOPC_burst_0_upstream_non_bursting_master_requests;
  wire             SS_OCT_SOPC_burst_0_upstream_read;
  wire    [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata_from_sa;
  wire             SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa;
  reg              SS_OCT_SOPC_burst_0_upstream_reg_firsttransfer;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_selected_burstcount;
  reg              SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable;
  wire             SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable2;
  wire             SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_transaction_burst_count;
  wire             SS_OCT_SOPC_burst_0_upstream_unreg_firsttransfer;
  wire             SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;
  wire             SS_OCT_SOPC_burst_0_upstream_waits_for_read;
  wire             SS_OCT_SOPC_burst_0_upstream_waits_for_write;
  wire             SS_OCT_SOPC_burst_0_upstream_write;
  wire    [255: 0] SS_OCT_SOPC_burst_0_upstream_writedata;
  wire             clock_crossing_master_ddr2_m1_arbiterlock;
  wire             clock_crossing_master_ddr2_m1_arbiterlock2;
  wire             clock_crossing_master_ddr2_m1_continuerequest;
  wire             clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_rdv_fifo_empty_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_rdv_fifo_output_from_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register;
  wire             clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_saved_grant_SS_OCT_SOPC_burst_0_upstream;
  reg              d1_SS_OCT_SOPC_burst_0_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_SS_OCT_SOPC_burst_0_upstream_load_fifo;
  wire             wait_for_SS_OCT_SOPC_burst_0_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~SS_OCT_SOPC_burst_0_upstream_end_xfer;
    end


  assign SS_OCT_SOPC_burst_0_upstream_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream));
  //assign SS_OCT_SOPC_burst_0_upstream_readdata_from_sa = SS_OCT_SOPC_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_readdata_from_sa = SS_OCT_SOPC_burst_0_upstream_readdata;

  assign clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream = (1) & (clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write);
  //assign SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa = SS_OCT_SOPC_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa = SS_OCT_SOPC_burst_0_upstream_waitrequest;

  //assign SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa = SS_OCT_SOPC_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa = SS_OCT_SOPC_burst_0_upstream_readdatavalid;

  //SS_OCT_SOPC_burst_0_upstream_arb_share_counter set values, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_arb_share_set_values = (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream)? (((clock_crossing_master_ddr2_m1_write) ? clock_crossing_master_ddr2_m1_burstcount : 1)) :
    1;

  //SS_OCT_SOPC_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_non_bursting_master_requests = 0;

  //SS_OCT_SOPC_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_any_bursting_master_saved_grant = clock_crossing_master_ddr2_m1_saved_grant_SS_OCT_SOPC_burst_0_upstream;

  //SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value = SS_OCT_SOPC_burst_0_upstream_firsttransfer ? (SS_OCT_SOPC_burst_0_upstream_arb_share_set_values - 1) : |SS_OCT_SOPC_burst_0_upstream_arb_share_counter ? (SS_OCT_SOPC_burst_0_upstream_arb_share_counter - 1) : 0;

  //SS_OCT_SOPC_burst_0_upstream_allgrants all slave grants, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_allgrants = |SS_OCT_SOPC_burst_0_upstream_grant_vector;

  //SS_OCT_SOPC_burst_0_upstream_end_xfer assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_end_xfer = ~(SS_OCT_SOPC_burst_0_upstream_waits_for_read | SS_OCT_SOPC_burst_0_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream = SS_OCT_SOPC_burst_0_upstream_end_xfer & (~SS_OCT_SOPC_burst_0_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //SS_OCT_SOPC_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream & SS_OCT_SOPC_burst_0_upstream_allgrants) | (end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream & ~SS_OCT_SOPC_burst_0_upstream_non_bursting_master_requests);

  //SS_OCT_SOPC_burst_0_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_arb_share_counter <= 0;
      else if (SS_OCT_SOPC_burst_0_upstream_arb_counter_enable)
          SS_OCT_SOPC_burst_0_upstream_arb_share_counter <= SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value;
    end


  //SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable <= 0;
      else if ((|SS_OCT_SOPC_burst_0_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream) | (end_xfer_arb_share_counter_term_SS_OCT_SOPC_burst_0_upstream & ~SS_OCT_SOPC_burst_0_upstream_non_bursting_master_requests))
          SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable <= |SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value;
    end


  //clock_crossing_master_ddr2/m1 SS_OCT_SOPC_burst_0/upstream arbiterlock, which is an e_assign
  assign clock_crossing_master_ddr2_m1_arbiterlock = SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable & clock_crossing_master_ddr2_m1_continuerequest;

  //SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable2 = |SS_OCT_SOPC_burst_0_upstream_arb_share_counter_next_value;

  //clock_crossing_master_ddr2/m1 SS_OCT_SOPC_burst_0/upstream arbiterlock2, which is an e_assign
  assign clock_crossing_master_ddr2_m1_arbiterlock2 = SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable2 & clock_crossing_master_ddr2_m1_continuerequest;

  //SS_OCT_SOPC_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_any_continuerequest = 1;

  //clock_crossing_master_ddr2_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_master_ddr2_m1_continuerequest = 1;

  assign clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream = clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream & ~((clock_crossing_master_ddr2_m1_read & ((clock_crossing_master_ddr2_m1_latency_counter != 0) | (1 < clock_crossing_master_ddr2_m1_latency_counter))));
  //unique name for SS_OCT_SOPC_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_move_on_to_next_transaction = SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst & SS_OCT_SOPC_burst_0_upstream_load_fifo;

  //the currently selected burstcount for SS_OCT_SOPC_burst_0_upstream, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_selected_burstcount = (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream)? clock_crossing_master_ddr2_m1_burstcount :
    1;

  //burstcount_fifo_for_SS_OCT_SOPC_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_SS_OCT_SOPC_burst_0_upstream_module burstcount_fifo_for_SS_OCT_SOPC_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (SS_OCT_SOPC_burst_0_upstream_selected_burstcount),
      .data_out             (SS_OCT_SOPC_burst_0_upstream_transaction_burst_count),
      .empty                (SS_OCT_SOPC_burst_0_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read & SS_OCT_SOPC_burst_0_upstream_load_fifo & ~(SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst & SS_OCT_SOPC_burst_0_upstream_burstcount_fifo_empty))
    );

  //SS_OCT_SOPC_burst_0_upstream current burst minus one, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_current_burst_minus_one = SS_OCT_SOPC_burst_0_upstream_current_burst - 1;

  //what to load in current_burst, for SS_OCT_SOPC_burst_0_upstream, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_next_burst_count = (((in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read) & ~SS_OCT_SOPC_burst_0_upstream_load_fifo))? SS_OCT_SOPC_burst_0_upstream_selected_burstcount :
    ((in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read & SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst & SS_OCT_SOPC_burst_0_upstream_burstcount_fifo_empty))? SS_OCT_SOPC_burst_0_upstream_selected_burstcount :
    (SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst)? SS_OCT_SOPC_burst_0_upstream_transaction_burst_count :
    SS_OCT_SOPC_burst_0_upstream_current_burst_minus_one;

  //the current burst count for SS_OCT_SOPC_burst_0_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_current_burst <= 0;
      else if (SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa | (~SS_OCT_SOPC_burst_0_upstream_load_fifo & (in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read)))
          SS_OCT_SOPC_burst_0_upstream_current_burst <= SS_OCT_SOPC_burst_0_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_SS_OCT_SOPC_burst_0_upstream_load_fifo = (~SS_OCT_SOPC_burst_0_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read) & SS_OCT_SOPC_burst_0_upstream_load_fifo))? 1 :
    ~SS_OCT_SOPC_burst_0_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read) & ~SS_OCT_SOPC_burst_0_upstream_load_fifo | SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst)
          SS_OCT_SOPC_burst_0_upstream_load_fifo <= p0_SS_OCT_SOPC_burst_0_upstream_load_fifo;
    end


  //the last cycle in the burst for SS_OCT_SOPC_burst_0_upstream, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_this_cycle_is_the_last_burst = ~(|SS_OCT_SOPC_burst_0_upstream_current_burst_minus_one) & SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_clock_crossing_master_ddr2_m1_to_SS_OCT_SOPC_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_clock_crossing_master_ddr2_m1_to_SS_OCT_SOPC_burst_0_upstream_module rdv_fifo_for_clock_crossing_master_ddr2_m1_to_SS_OCT_SOPC_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream),
      .data_out             (clock_crossing_master_ddr2_m1_rdv_fifo_output_from_SS_OCT_SOPC_burst_0_upstream),
      .empty                (),
      .fifo_contains_ones_n (clock_crossing_master_ddr2_m1_rdv_fifo_empty_SS_OCT_SOPC_burst_0_upstream),
      .full                 (),
      .read                 (SS_OCT_SOPC_burst_0_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~SS_OCT_SOPC_burst_0_upstream_waits_for_read)
    );

  assign clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register = ~clock_crossing_master_ddr2_m1_rdv_fifo_empty_SS_OCT_SOPC_burst_0_upstream;
  //local readdatavalid clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream, which is an e_mux
  assign clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream = SS_OCT_SOPC_burst_0_upstream_readdatavalid_from_sa;

  //SS_OCT_SOPC_burst_0_upstream_writedata mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_writedata = clock_crossing_master_ddr2_m1_writedata;

  //byteaddress mux for SS_OCT_SOPC_burst_0/upstream, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_byteaddress = clock_crossing_master_ddr2_m1_address_to_slave;

  //master is always granted when requested
  assign clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream = clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream;

  //clock_crossing_master_ddr2/m1 saved-grant SS_OCT_SOPC_burst_0/upstream, which is an e_assign
  assign clock_crossing_master_ddr2_m1_saved_grant_SS_OCT_SOPC_burst_0_upstream = clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream;

  //allow new arb cycle for SS_OCT_SOPC_burst_0/upstream, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign SS_OCT_SOPC_burst_0_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign SS_OCT_SOPC_burst_0_upstream_master_qreq_vector = 1;

  //SS_OCT_SOPC_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_firsttransfer = SS_OCT_SOPC_burst_0_upstream_begins_xfer ? SS_OCT_SOPC_burst_0_upstream_unreg_firsttransfer : SS_OCT_SOPC_burst_0_upstream_reg_firsttransfer;

  //SS_OCT_SOPC_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_unreg_firsttransfer = ~(SS_OCT_SOPC_burst_0_upstream_slavearbiterlockenable & SS_OCT_SOPC_burst_0_upstream_any_continuerequest);

  //SS_OCT_SOPC_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_reg_firsttransfer <= 1'b1;
      else if (SS_OCT_SOPC_burst_0_upstream_begins_xfer)
          SS_OCT_SOPC_burst_0_upstream_reg_firsttransfer <= SS_OCT_SOPC_burst_0_upstream_unreg_firsttransfer;
    end


  //SS_OCT_SOPC_burst_0_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_next_bbt_burstcount = ((((SS_OCT_SOPC_burst_0_upstream_write) && (SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter == 0))))? (SS_OCT_SOPC_burst_0_upstream_burstcount - 1) :
    ((((SS_OCT_SOPC_burst_0_upstream_read) && (SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter == 0))))? 0 :
    (SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter - 1);

  //SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter <= 0;
      else if (SS_OCT_SOPC_burst_0_upstream_begins_xfer)
          SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter <= SS_OCT_SOPC_burst_0_upstream_next_bbt_burstcount;
    end


  //SS_OCT_SOPC_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_beginbursttransfer_internal = SS_OCT_SOPC_burst_0_upstream_begins_xfer & (SS_OCT_SOPC_burst_0_upstream_bbt_burstcounter == 0);

  //SS_OCT_SOPC_burst_0_upstream_read assignment, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_read = clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream & clock_crossing_master_ddr2_m1_read;

  //SS_OCT_SOPC_burst_0_upstream_write assignment, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_write = clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream & clock_crossing_master_ddr2_m1_write;

  //SS_OCT_SOPC_burst_0_upstream_address mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_address = clock_crossing_master_ddr2_m1_address_to_slave;

  //d1_SS_OCT_SOPC_burst_0_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_SS_OCT_SOPC_burst_0_upstream_end_xfer <= 1;
      else 
        d1_SS_OCT_SOPC_burst_0_upstream_end_xfer <= SS_OCT_SOPC_burst_0_upstream_end_xfer;
    end


  //SS_OCT_SOPC_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_waits_for_read = SS_OCT_SOPC_burst_0_upstream_in_a_read_cycle & SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;

  //SS_OCT_SOPC_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_in_a_read_cycle = clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream & clock_crossing_master_ddr2_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = SS_OCT_SOPC_burst_0_upstream_in_a_read_cycle;

  //SS_OCT_SOPC_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_waits_for_write = SS_OCT_SOPC_burst_0_upstream_in_a_write_cycle & SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;

  //SS_OCT_SOPC_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_upstream_in_a_write_cycle = clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream & clock_crossing_master_ddr2_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = SS_OCT_SOPC_burst_0_upstream_in_a_write_cycle;

  assign wait_for_SS_OCT_SOPC_burst_0_upstream_counter = 0;
  //SS_OCT_SOPC_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_byteenable = (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream)? clock_crossing_master_ddr2_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_burstcount = (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream)? clock_crossing_master_ddr2_m1_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //SS_OCT_SOPC_burst_0/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //clock_crossing_master_ddr2/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream && (clock_crossing_master_ddr2_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: clock_crossing_master_ddr2/m1 drove 0 on its 'burstcount' port while accessing slave SS_OCT_SOPC_burst_0/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_burst_0_downstream_arbitrator (
                                                   // inputs:
                                                    SS_OCT_SOPC_burst_0_downstream_address,
                                                    SS_OCT_SOPC_burst_0_downstream_burstcount,
                                                    SS_OCT_SOPC_burst_0_downstream_byteenable,
                                                    SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1,
                                                    SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1,
                                                    SS_OCT_SOPC_burst_0_downstream_read,
                                                    SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1,
                                                    SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register,
                                                    SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1,
                                                    SS_OCT_SOPC_burst_0_downstream_write,
                                                    SS_OCT_SOPC_burst_0_downstream_writedata,
                                                    clk,
                                                    d1_ddr2_s1_end_xfer,
                                                    ddr2_s1_readdata_from_sa,
                                                    ddr2_s1_waitrequest_n_from_sa,
                                                    reset_n,

                                                   // outputs:
                                                    SS_OCT_SOPC_burst_0_downstream_address_to_slave,
                                                    SS_OCT_SOPC_burst_0_downstream_latency_counter,
                                                    SS_OCT_SOPC_burst_0_downstream_readdata,
                                                    SS_OCT_SOPC_burst_0_downstream_readdatavalid,
                                                    SS_OCT_SOPC_burst_0_downstream_reset_n,
                                                    SS_OCT_SOPC_burst_0_downstream_waitrequest
                                                 )
;

  output  [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address_to_slave;
  output           SS_OCT_SOPC_burst_0_downstream_latency_counter;
  output  [255: 0] SS_OCT_SOPC_burst_0_downstream_readdata;
  output           SS_OCT_SOPC_burst_0_downstream_readdatavalid;
  output           SS_OCT_SOPC_burst_0_downstream_reset_n;
  output           SS_OCT_SOPC_burst_0_downstream_waitrequest;
  input   [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address;
  input   [  2: 0] SS_OCT_SOPC_burst_0_downstream_burstcount;
  input   [ 31: 0] SS_OCT_SOPC_burst_0_downstream_byteenable;
  input            SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1;
  input            SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1;
  input            SS_OCT_SOPC_burst_0_downstream_read;
  input            SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1;
  input            SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register;
  input            SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1;
  input            SS_OCT_SOPC_burst_0_downstream_write;
  input   [255: 0] SS_OCT_SOPC_burst_0_downstream_writedata;
  input            clk;
  input            d1_ddr2_s1_end_xfer;
  input   [255: 0] ddr2_s1_readdata_from_sa;
  input            ddr2_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg     [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address_last_time;
  wire    [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address_to_slave;
  reg     [  2: 0] SS_OCT_SOPC_burst_0_downstream_burstcount_last_time;
  reg     [ 31: 0] SS_OCT_SOPC_burst_0_downstream_byteenable_last_time;
  wire             SS_OCT_SOPC_burst_0_downstream_is_granted_some_slave;
  reg              SS_OCT_SOPC_burst_0_downstream_latency_counter;
  reg              SS_OCT_SOPC_burst_0_downstream_read_but_no_slave_selected;
  reg              SS_OCT_SOPC_burst_0_downstream_read_last_time;
  wire    [255: 0] SS_OCT_SOPC_burst_0_downstream_readdata;
  wire             SS_OCT_SOPC_burst_0_downstream_readdatavalid;
  wire             SS_OCT_SOPC_burst_0_downstream_reset_n;
  wire             SS_OCT_SOPC_burst_0_downstream_run;
  wire             SS_OCT_SOPC_burst_0_downstream_waitrequest;
  reg              SS_OCT_SOPC_burst_0_downstream_write_last_time;
  reg     [255: 0] SS_OCT_SOPC_burst_0_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_SS_OCT_SOPC_burst_0_downstream_latency_counter;
  wire             pre_flush_SS_OCT_SOPC_burst_0_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1 | ~SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1) & (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 | ~SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1) & ((~SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1 | ~(SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write) | (1 & ddr2_s1_waitrequest_n_from_sa & (SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write)))) & ((~SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1 | ~(SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write) | (1 & ddr2_s1_waitrequest_n_from_sa & (SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign SS_OCT_SOPC_burst_0_downstream_address_to_slave = SS_OCT_SOPC_burst_0_downstream_address;

  //SS_OCT_SOPC_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_read_but_no_slave_selected <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_read_but_no_slave_selected <= SS_OCT_SOPC_burst_0_downstream_read & SS_OCT_SOPC_burst_0_downstream_run & ~SS_OCT_SOPC_burst_0_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign SS_OCT_SOPC_burst_0_downstream_is_granted_some_slave = SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_SS_OCT_SOPC_burst_0_downstream_readdatavalid = SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign SS_OCT_SOPC_burst_0_downstream_readdatavalid = SS_OCT_SOPC_burst_0_downstream_read_but_no_slave_selected |
    pre_flush_SS_OCT_SOPC_burst_0_downstream_readdatavalid;

  //SS_OCT_SOPC_burst_0/downstream readdata mux, which is an e_mux
  assign SS_OCT_SOPC_burst_0_downstream_readdata = ddr2_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_waitrequest = ~SS_OCT_SOPC_burst_0_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_latency_counter <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_latency_counter <= p1_SS_OCT_SOPC_burst_0_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_SS_OCT_SOPC_burst_0_downstream_latency_counter = ((SS_OCT_SOPC_burst_0_downstream_run & SS_OCT_SOPC_burst_0_downstream_read))? latency_load_value :
    (SS_OCT_SOPC_burst_0_downstream_latency_counter)? SS_OCT_SOPC_burst_0_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //SS_OCT_SOPC_burst_0_downstream_reset_n assignment, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //SS_OCT_SOPC_burst_0_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_address_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_address_last_time <= SS_OCT_SOPC_burst_0_downstream_address;
    end


  //SS_OCT_SOPC_burst_0/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= SS_OCT_SOPC_burst_0_downstream_waitrequest & (SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write);
    end


  //SS_OCT_SOPC_burst_0_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_address != SS_OCT_SOPC_burst_0_downstream_address_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_burstcount_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_burstcount_last_time <= SS_OCT_SOPC_burst_0_downstream_burstcount;
    end


  //SS_OCT_SOPC_burst_0_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_burstcount != SS_OCT_SOPC_burst_0_downstream_burstcount_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_byteenable_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_byteenable_last_time <= SS_OCT_SOPC_burst_0_downstream_byteenable;
    end


  //SS_OCT_SOPC_burst_0_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_byteenable != SS_OCT_SOPC_burst_0_downstream_byteenable_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_read_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_read_last_time <= SS_OCT_SOPC_burst_0_downstream_read;
    end


  //SS_OCT_SOPC_burst_0_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_read != SS_OCT_SOPC_burst_0_downstream_read_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_write_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_write_last_time <= SS_OCT_SOPC_burst_0_downstream_write;
    end


  //SS_OCT_SOPC_burst_0_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_write != SS_OCT_SOPC_burst_0_downstream_write_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_burst_0_downstream_writedata_last_time <= 0;
      else 
        SS_OCT_SOPC_burst_0_downstream_writedata_last_time <= SS_OCT_SOPC_burst_0_downstream_writedata;
    end


  //SS_OCT_SOPC_burst_0_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_burst_0_downstream_writedata != SS_OCT_SOPC_burst_0_downstream_writedata_last_time) & SS_OCT_SOPC_burst_0_downstream_write)
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_clock_0_in_arbitrator (
                                           // inputs:
                                            SS_OCT_SOPC_clock_0_in_endofpacket,
                                            SS_OCT_SOPC_clock_0_in_readdata,
                                            SS_OCT_SOPC_clock_0_in_waitrequest,
                                            clk,
                                            cpu_data_master_address_to_slave,
                                            cpu_data_master_byteenable,
                                            cpu_data_master_latency_counter,
                                            cpu_data_master_read,
                                            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                            cpu_data_master_write,
                                            cpu_data_master_writedata,
                                            reset_n,

                                           // outputs:
                                            SS_OCT_SOPC_clock_0_in_address,
                                            SS_OCT_SOPC_clock_0_in_byteenable,
                                            SS_OCT_SOPC_clock_0_in_endofpacket_from_sa,
                                            SS_OCT_SOPC_clock_0_in_nativeaddress,
                                            SS_OCT_SOPC_clock_0_in_read,
                                            SS_OCT_SOPC_clock_0_in_readdata_from_sa,
                                            SS_OCT_SOPC_clock_0_in_reset_n,
                                            SS_OCT_SOPC_clock_0_in_waitrequest_from_sa,
                                            SS_OCT_SOPC_clock_0_in_write,
                                            SS_OCT_SOPC_clock_0_in_writedata,
                                            cpu_data_master_granted_SS_OCT_SOPC_clock_0_in,
                                            cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in,
                                            cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in,
                                            cpu_data_master_requests_SS_OCT_SOPC_clock_0_in,
                                            d1_SS_OCT_SOPC_clock_0_in_end_xfer
                                         )
;

  output  [  3: 0] SS_OCT_SOPC_clock_0_in_address;
  output  [  1: 0] SS_OCT_SOPC_clock_0_in_byteenable;
  output           SS_OCT_SOPC_clock_0_in_endofpacket_from_sa;
  output  [  2: 0] SS_OCT_SOPC_clock_0_in_nativeaddress;
  output           SS_OCT_SOPC_clock_0_in_read;
  output  [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata_from_sa;
  output           SS_OCT_SOPC_clock_0_in_reset_n;
  output           SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;
  output           SS_OCT_SOPC_clock_0_in_write;
  output  [ 15: 0] SS_OCT_SOPC_clock_0_in_writedata;
  output           cpu_data_master_granted_SS_OCT_SOPC_clock_0_in;
  output           cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in;
  output           cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in;
  output           cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;
  output           d1_SS_OCT_SOPC_clock_0_in_end_xfer;
  input            SS_OCT_SOPC_clock_0_in_endofpacket;
  input   [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata;
  input            SS_OCT_SOPC_clock_0_in_waitrequest;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] SS_OCT_SOPC_clock_0_in_address;
  wire             SS_OCT_SOPC_clock_0_in_allgrants;
  wire             SS_OCT_SOPC_clock_0_in_allow_new_arb_cycle;
  wire             SS_OCT_SOPC_clock_0_in_any_bursting_master_saved_grant;
  wire             SS_OCT_SOPC_clock_0_in_any_continuerequest;
  wire             SS_OCT_SOPC_clock_0_in_arb_counter_enable;
  reg     [  1: 0] SS_OCT_SOPC_clock_0_in_arb_share_counter;
  wire    [  1: 0] SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value;
  wire    [  1: 0] SS_OCT_SOPC_clock_0_in_arb_share_set_values;
  wire             SS_OCT_SOPC_clock_0_in_beginbursttransfer_internal;
  wire             SS_OCT_SOPC_clock_0_in_begins_xfer;
  wire    [  1: 0] SS_OCT_SOPC_clock_0_in_byteenable;
  wire             SS_OCT_SOPC_clock_0_in_end_xfer;
  wire             SS_OCT_SOPC_clock_0_in_endofpacket_from_sa;
  wire             SS_OCT_SOPC_clock_0_in_firsttransfer;
  wire             SS_OCT_SOPC_clock_0_in_grant_vector;
  wire             SS_OCT_SOPC_clock_0_in_in_a_read_cycle;
  wire             SS_OCT_SOPC_clock_0_in_in_a_write_cycle;
  wire             SS_OCT_SOPC_clock_0_in_master_qreq_vector;
  wire    [  2: 0] SS_OCT_SOPC_clock_0_in_nativeaddress;
  wire             SS_OCT_SOPC_clock_0_in_non_bursting_master_requests;
  wire             SS_OCT_SOPC_clock_0_in_read;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata_from_sa;
  reg              SS_OCT_SOPC_clock_0_in_reg_firsttransfer;
  wire             SS_OCT_SOPC_clock_0_in_reset_n;
  reg              SS_OCT_SOPC_clock_0_in_slavearbiterlockenable;
  wire             SS_OCT_SOPC_clock_0_in_slavearbiterlockenable2;
  wire             SS_OCT_SOPC_clock_0_in_unreg_firsttransfer;
  wire             SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;
  wire             SS_OCT_SOPC_clock_0_in_waits_for_read;
  wire             SS_OCT_SOPC_clock_0_in_waits_for_write;
  wire             SS_OCT_SOPC_clock_0_in_write;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_in_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_saved_grant_SS_OCT_SOPC_clock_0_in;
  reg              d1_SS_OCT_SOPC_clock_0_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_SS_OCT_SOPC_clock_0_in_from_cpu_data_master;
  wire             wait_for_SS_OCT_SOPC_clock_0_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~SS_OCT_SOPC_clock_0_in_end_xfer;
    end


  assign SS_OCT_SOPC_clock_0_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in));
  //assign SS_OCT_SOPC_clock_0_in_readdata_from_sa = SS_OCT_SOPC_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_readdata_from_sa = SS_OCT_SOPC_clock_0_in_readdata;

  assign cpu_data_master_requests_SS_OCT_SOPC_clock_0_in = ({cpu_data_master_address_to_slave[30 : 5] , 5'b0} == 31'h48112400) & (cpu_data_master_read | cpu_data_master_write);
  //assign SS_OCT_SOPC_clock_0_in_waitrequest_from_sa = SS_OCT_SOPC_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_waitrequest_from_sa = SS_OCT_SOPC_clock_0_in_waitrequest;

  //SS_OCT_SOPC_clock_0_in_arb_share_counter set values, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_arb_share_set_values = 1;

  //SS_OCT_SOPC_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_non_bursting_master_requests = cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;

  //SS_OCT_SOPC_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_any_bursting_master_saved_grant = 0;

  //SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value = SS_OCT_SOPC_clock_0_in_firsttransfer ? (SS_OCT_SOPC_clock_0_in_arb_share_set_values - 1) : |SS_OCT_SOPC_clock_0_in_arb_share_counter ? (SS_OCT_SOPC_clock_0_in_arb_share_counter - 1) : 0;

  //SS_OCT_SOPC_clock_0_in_allgrants all slave grants, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_allgrants = |SS_OCT_SOPC_clock_0_in_grant_vector;

  //SS_OCT_SOPC_clock_0_in_end_xfer assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_end_xfer = ~(SS_OCT_SOPC_clock_0_in_waits_for_read | SS_OCT_SOPC_clock_0_in_waits_for_write);

  //end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in = SS_OCT_SOPC_clock_0_in_end_xfer & (~SS_OCT_SOPC_clock_0_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //SS_OCT_SOPC_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_arb_counter_enable = (end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in & SS_OCT_SOPC_clock_0_in_allgrants) | (end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in & ~SS_OCT_SOPC_clock_0_in_non_bursting_master_requests);

  //SS_OCT_SOPC_clock_0_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_in_arb_share_counter <= 0;
      else if (SS_OCT_SOPC_clock_0_in_arb_counter_enable)
          SS_OCT_SOPC_clock_0_in_arb_share_counter <= SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value;
    end


  //SS_OCT_SOPC_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_in_slavearbiterlockenable <= 0;
      else if ((|SS_OCT_SOPC_clock_0_in_master_qreq_vector & end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in) | (end_xfer_arb_share_counter_term_SS_OCT_SOPC_clock_0_in & ~SS_OCT_SOPC_clock_0_in_non_bursting_master_requests))
          SS_OCT_SOPC_clock_0_in_slavearbiterlockenable <= |SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value;
    end


  //cpu/data_master SS_OCT_SOPC_clock_0/in arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = SS_OCT_SOPC_clock_0_in_slavearbiterlockenable & cpu_data_master_continuerequest;

  //SS_OCT_SOPC_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_slavearbiterlockenable2 = |SS_OCT_SOPC_clock_0_in_arb_share_counter_next_value;

  //cpu/data_master SS_OCT_SOPC_clock_0/in arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = SS_OCT_SOPC_clock_0_in_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //SS_OCT_SOPC_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in = cpu_data_master_requests_SS_OCT_SOPC_clock_0_in & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in, which is an e_mux
  assign cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in & cpu_data_master_read & ~SS_OCT_SOPC_clock_0_in_waits_for_read;

  //SS_OCT_SOPC_clock_0_in_writedata mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_writedata = cpu_data_master_writedata;

  //assign SS_OCT_SOPC_clock_0_in_endofpacket_from_sa = SS_OCT_SOPC_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_endofpacket_from_sa = SS_OCT_SOPC_clock_0_in_endofpacket;

  //master is always granted when requested
  assign cpu_data_master_granted_SS_OCT_SOPC_clock_0_in = cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in;

  //cpu/data_master saved-grant SS_OCT_SOPC_clock_0/in, which is an e_assign
  assign cpu_data_master_saved_grant_SS_OCT_SOPC_clock_0_in = cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;

  //allow new arb cycle for SS_OCT_SOPC_clock_0/in, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign SS_OCT_SOPC_clock_0_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign SS_OCT_SOPC_clock_0_in_master_qreq_vector = 1;

  //SS_OCT_SOPC_clock_0_in_reset_n assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_reset_n = reset_n;

  //SS_OCT_SOPC_clock_0_in_firsttransfer first transaction, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_firsttransfer = SS_OCT_SOPC_clock_0_in_begins_xfer ? SS_OCT_SOPC_clock_0_in_unreg_firsttransfer : SS_OCT_SOPC_clock_0_in_reg_firsttransfer;

  //SS_OCT_SOPC_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_unreg_firsttransfer = ~(SS_OCT_SOPC_clock_0_in_slavearbiterlockenable & SS_OCT_SOPC_clock_0_in_any_continuerequest);

  //SS_OCT_SOPC_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_in_reg_firsttransfer <= 1'b1;
      else if (SS_OCT_SOPC_clock_0_in_begins_xfer)
          SS_OCT_SOPC_clock_0_in_reg_firsttransfer <= SS_OCT_SOPC_clock_0_in_unreg_firsttransfer;
    end


  //SS_OCT_SOPC_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_beginbursttransfer_internal = SS_OCT_SOPC_clock_0_in_begins_xfer;

  //SS_OCT_SOPC_clock_0_in_read assignment, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_read = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in & cpu_data_master_read;

  //SS_OCT_SOPC_clock_0_in_write assignment, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_write = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in & cpu_data_master_write;

  assign shifted_address_to_SS_OCT_SOPC_clock_0_in_from_cpu_data_master = cpu_data_master_address_to_slave;
  //SS_OCT_SOPC_clock_0_in_address mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_address = shifted_address_to_SS_OCT_SOPC_clock_0_in_from_cpu_data_master >> 2;

  //slaveid SS_OCT_SOPC_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_nativeaddress = cpu_data_master_address_to_slave >> 2;

  //d1_SS_OCT_SOPC_clock_0_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_SS_OCT_SOPC_clock_0_in_end_xfer <= 1;
      else 
        d1_SS_OCT_SOPC_clock_0_in_end_xfer <= SS_OCT_SOPC_clock_0_in_end_xfer;
    end


  //SS_OCT_SOPC_clock_0_in_waits_for_read in a cycle, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_waits_for_read = SS_OCT_SOPC_clock_0_in_in_a_read_cycle & SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;

  //SS_OCT_SOPC_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_in_a_read_cycle = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = SS_OCT_SOPC_clock_0_in_in_a_read_cycle;

  //SS_OCT_SOPC_clock_0_in_waits_for_write in a cycle, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_waits_for_write = SS_OCT_SOPC_clock_0_in_in_a_write_cycle & SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;

  //SS_OCT_SOPC_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_in_in_a_write_cycle = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = SS_OCT_SOPC_clock_0_in_in_a_write_cycle;

  assign wait_for_SS_OCT_SOPC_clock_0_in_counter = 0;
  //SS_OCT_SOPC_clock_0_in_byteenable byte enable port mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_in_byteenable = (cpu_data_master_granted_SS_OCT_SOPC_clock_0_in)? cpu_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //SS_OCT_SOPC_clock_0/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_clock_0_out_arbitrator (
                                            // inputs:
                                             SS_OCT_SOPC_clock_0_out_address,
                                             SS_OCT_SOPC_clock_0_out_byteenable,
                                             SS_OCT_SOPC_clock_0_out_granted_pll_s1,
                                             SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1,
                                             SS_OCT_SOPC_clock_0_out_read,
                                             SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1,
                                             SS_OCT_SOPC_clock_0_out_requests_pll_s1,
                                             SS_OCT_SOPC_clock_0_out_write,
                                             SS_OCT_SOPC_clock_0_out_writedata,
                                             clk,
                                             d1_pll_s1_end_xfer,
                                             pll_s1_readdata_from_sa,
                                             reset_n,

                                            // outputs:
                                             SS_OCT_SOPC_clock_0_out_address_to_slave,
                                             SS_OCT_SOPC_clock_0_out_readdata,
                                             SS_OCT_SOPC_clock_0_out_reset_n,
                                             SS_OCT_SOPC_clock_0_out_waitrequest
                                          )
;

  output  [  3: 0] SS_OCT_SOPC_clock_0_out_address_to_slave;
  output  [ 15: 0] SS_OCT_SOPC_clock_0_out_readdata;
  output           SS_OCT_SOPC_clock_0_out_reset_n;
  output           SS_OCT_SOPC_clock_0_out_waitrequest;
  input   [  3: 0] SS_OCT_SOPC_clock_0_out_address;
  input   [  1: 0] SS_OCT_SOPC_clock_0_out_byteenable;
  input            SS_OCT_SOPC_clock_0_out_granted_pll_s1;
  input            SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1;
  input            SS_OCT_SOPC_clock_0_out_read;
  input            SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1;
  input            SS_OCT_SOPC_clock_0_out_requests_pll_s1;
  input            SS_OCT_SOPC_clock_0_out_write;
  input   [ 15: 0] SS_OCT_SOPC_clock_0_out_writedata;
  input            clk;
  input            d1_pll_s1_end_xfer;
  input   [ 15: 0] pll_s1_readdata_from_sa;
  input            reset_n;

  reg     [  3: 0] SS_OCT_SOPC_clock_0_out_address_last_time;
  wire    [  3: 0] SS_OCT_SOPC_clock_0_out_address_to_slave;
  reg     [  1: 0] SS_OCT_SOPC_clock_0_out_byteenable_last_time;
  reg              SS_OCT_SOPC_clock_0_out_read_last_time;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_out_readdata;
  wire             SS_OCT_SOPC_clock_0_out_reset_n;
  wire             SS_OCT_SOPC_clock_0_out_run;
  wire             SS_OCT_SOPC_clock_0_out_waitrequest;
  reg              SS_OCT_SOPC_clock_0_out_write_last_time;
  reg     [ 15: 0] SS_OCT_SOPC_clock_0_out_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             r_2;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & ((~SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1 | ~SS_OCT_SOPC_clock_0_out_read | (1 & ~d1_pll_s1_end_xfer & SS_OCT_SOPC_clock_0_out_read))) & ((~SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1 | ~SS_OCT_SOPC_clock_0_out_write | (1 & SS_OCT_SOPC_clock_0_out_write)));

  //cascaded wait assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign SS_OCT_SOPC_clock_0_out_address_to_slave = SS_OCT_SOPC_clock_0_out_address;

  //SS_OCT_SOPC_clock_0/out readdata mux, which is an e_mux
  assign SS_OCT_SOPC_clock_0_out_readdata = pll_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_waitrequest = ~SS_OCT_SOPC_clock_0_out_run;

  //SS_OCT_SOPC_clock_0_out_reset_n assignment, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //SS_OCT_SOPC_clock_0_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_out_address_last_time <= 0;
      else 
        SS_OCT_SOPC_clock_0_out_address_last_time <= SS_OCT_SOPC_clock_0_out_address;
    end


  //SS_OCT_SOPC_clock_0/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= SS_OCT_SOPC_clock_0_out_waitrequest & (SS_OCT_SOPC_clock_0_out_read | SS_OCT_SOPC_clock_0_out_write);
    end


  //SS_OCT_SOPC_clock_0_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_clock_0_out_address != SS_OCT_SOPC_clock_0_out_address_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_clock_0_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_clock_0_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_out_byteenable_last_time <= 0;
      else 
        SS_OCT_SOPC_clock_0_out_byteenable_last_time <= SS_OCT_SOPC_clock_0_out_byteenable;
    end


  //SS_OCT_SOPC_clock_0_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_clock_0_out_byteenable != SS_OCT_SOPC_clock_0_out_byteenable_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_clock_0_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_clock_0_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_out_read_last_time <= 0;
      else 
        SS_OCT_SOPC_clock_0_out_read_last_time <= SS_OCT_SOPC_clock_0_out_read;
    end


  //SS_OCT_SOPC_clock_0_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_clock_0_out_read != SS_OCT_SOPC_clock_0_out_read_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_clock_0_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_clock_0_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_out_write_last_time <= 0;
      else 
        SS_OCT_SOPC_clock_0_out_write_last_time <= SS_OCT_SOPC_clock_0_out_write;
    end


  //SS_OCT_SOPC_clock_0_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_clock_0_out_write != SS_OCT_SOPC_clock_0_out_write_last_time))
        begin
          $write("%0d ns: SS_OCT_SOPC_clock_0_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_clock_0_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          SS_OCT_SOPC_clock_0_out_writedata_last_time <= 0;
      else 
        SS_OCT_SOPC_clock_0_out_writedata_last_time <= SS_OCT_SOPC_clock_0_out_writedata;
    end


  //SS_OCT_SOPC_clock_0_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (SS_OCT_SOPC_clock_0_out_writedata != SS_OCT_SOPC_clock_0_out_writedata_last_time) & SS_OCT_SOPC_clock_0_out_write)
        begin
          $write("%0d ns: SS_OCT_SOPC_clock_0_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_clock_crossing_ddr2_cpu_s1_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p96_full_96;
  wire             p96_stage_96;
  wire             p97_full_97;
  wire             p97_stage_97;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  reg              stage_96;
  reg              stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_ddr2_cpu_s1_arbitrator (
                                               // inputs:
                                                clk,
                                                clock_crossing_ddr2_cpu_s1_endofpacket,
                                                clock_crossing_ddr2_cpu_s1_readdata,
                                                clock_crossing_ddr2_cpu_s1_readdatavalid,
                                                clock_crossing_ddr2_cpu_s1_waitrequest,
                                                cpu_data_master_address_to_slave,
                                                cpu_data_master_byteenable,
                                                cpu_data_master_latency_counter,
                                                cpu_data_master_read,
                                                cpu_data_master_write,
                                                cpu_data_master_writedata,
                                                reset_n,

                                               // outputs:
                                                clock_crossing_ddr2_cpu_s1_address,
                                                clock_crossing_ddr2_cpu_s1_byteenable,
                                                clock_crossing_ddr2_cpu_s1_endofpacket_from_sa,
                                                clock_crossing_ddr2_cpu_s1_nativeaddress,
                                                clock_crossing_ddr2_cpu_s1_read,
                                                clock_crossing_ddr2_cpu_s1_readdata_from_sa,
                                                clock_crossing_ddr2_cpu_s1_reset_n,
                                                clock_crossing_ddr2_cpu_s1_waitrequest_from_sa,
                                                clock_crossing_ddr2_cpu_s1_write,
                                                clock_crossing_ddr2_cpu_s1_writedata,
                                                cpu_data_master_granted_clock_crossing_ddr2_cpu_s1,
                                                cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1,
                                                cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1,
                                                cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                                cpu_data_master_requests_clock_crossing_ddr2_cpu_s1,
                                                d1_clock_crossing_ddr2_cpu_s1_end_xfer
                                             )
;

  output  [ 27: 0] clock_crossing_ddr2_cpu_s1_address;
  output  [  3: 0] clock_crossing_ddr2_cpu_s1_byteenable;
  output           clock_crossing_ddr2_cpu_s1_endofpacket_from_sa;
  output  [ 27: 0] clock_crossing_ddr2_cpu_s1_nativeaddress;
  output           clock_crossing_ddr2_cpu_s1_read;
  output  [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata_from_sa;
  output           clock_crossing_ddr2_cpu_s1_reset_n;
  output           clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;
  output           clock_crossing_ddr2_cpu_s1_write;
  output  [ 31: 0] clock_crossing_ddr2_cpu_s1_writedata;
  output           cpu_data_master_granted_clock_crossing_ddr2_cpu_s1;
  output           cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1;
  output           cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1;
  output           cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  output           cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;
  output           d1_clock_crossing_ddr2_cpu_s1_end_xfer;
  input            clk;
  input            clock_crossing_ddr2_cpu_s1_endofpacket;
  input   [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata;
  input            clock_crossing_ddr2_cpu_s1_readdatavalid;
  input            clock_crossing_ddr2_cpu_s1_waitrequest;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [ 27: 0] clock_crossing_ddr2_cpu_s1_address;
  wire             clock_crossing_ddr2_cpu_s1_allgrants;
  wire             clock_crossing_ddr2_cpu_s1_allow_new_arb_cycle;
  wire             clock_crossing_ddr2_cpu_s1_any_bursting_master_saved_grant;
  wire             clock_crossing_ddr2_cpu_s1_any_continuerequest;
  wire             clock_crossing_ddr2_cpu_s1_arb_counter_enable;
  reg     [  1: 0] clock_crossing_ddr2_cpu_s1_arb_share_counter;
  wire    [  1: 0] clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value;
  wire    [  1: 0] clock_crossing_ddr2_cpu_s1_arb_share_set_values;
  wire             clock_crossing_ddr2_cpu_s1_beginbursttransfer_internal;
  wire             clock_crossing_ddr2_cpu_s1_begins_xfer;
  wire    [  3: 0] clock_crossing_ddr2_cpu_s1_byteenable;
  wire             clock_crossing_ddr2_cpu_s1_end_xfer;
  wire             clock_crossing_ddr2_cpu_s1_endofpacket_from_sa;
  wire             clock_crossing_ddr2_cpu_s1_firsttransfer;
  wire             clock_crossing_ddr2_cpu_s1_grant_vector;
  wire             clock_crossing_ddr2_cpu_s1_in_a_read_cycle;
  wire             clock_crossing_ddr2_cpu_s1_in_a_write_cycle;
  wire             clock_crossing_ddr2_cpu_s1_master_qreq_vector;
  wire             clock_crossing_ddr2_cpu_s1_move_on_to_next_transaction;
  wire    [ 27: 0] clock_crossing_ddr2_cpu_s1_nativeaddress;
  wire             clock_crossing_ddr2_cpu_s1_non_bursting_master_requests;
  wire             clock_crossing_ddr2_cpu_s1_read;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata_from_sa;
  wire             clock_crossing_ddr2_cpu_s1_readdatavalid_from_sa;
  reg              clock_crossing_ddr2_cpu_s1_reg_firsttransfer;
  wire             clock_crossing_ddr2_cpu_s1_reset_n;
  reg              clock_crossing_ddr2_cpu_s1_slavearbiterlockenable;
  wire             clock_crossing_ddr2_cpu_s1_slavearbiterlockenable2;
  wire             clock_crossing_ddr2_cpu_s1_unreg_firsttransfer;
  wire             clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;
  wire             clock_crossing_ddr2_cpu_s1_waits_for_read;
  wire             clock_crossing_ddr2_cpu_s1_waits_for_write;
  wire             clock_crossing_ddr2_cpu_s1_write;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_s1_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_rdv_fifo_empty_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_rdv_fifo_output_from_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  wire             cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_saved_grant_clock_crossing_ddr2_cpu_s1;
  reg              d1_clock_crossing_ddr2_cpu_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_clock_crossing_ddr2_cpu_s1_from_cpu_data_master;
  wire             wait_for_clock_crossing_ddr2_cpu_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~clock_crossing_ddr2_cpu_s1_end_xfer;
    end


  assign clock_crossing_ddr2_cpu_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1));
  //assign clock_crossing_ddr2_cpu_s1_readdatavalid_from_sa = clock_crossing_ddr2_cpu_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_readdatavalid_from_sa = clock_crossing_ddr2_cpu_s1_readdatavalid;

  //assign clock_crossing_ddr2_cpu_s1_readdata_from_sa = clock_crossing_ddr2_cpu_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_readdata_from_sa = clock_crossing_ddr2_cpu_s1_readdata;

  assign cpu_data_master_requests_clock_crossing_ddr2_cpu_s1 = ({cpu_data_master_address_to_slave[30] , 30'b0} == 31'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign clock_crossing_ddr2_cpu_s1_waitrequest_from_sa = clock_crossing_ddr2_cpu_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_waitrequest_from_sa = clock_crossing_ddr2_cpu_s1_waitrequest;

  //clock_crossing_ddr2_cpu_s1_arb_share_counter set values, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_arb_share_set_values = 1;

  //clock_crossing_ddr2_cpu_s1_non_bursting_master_requests mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_non_bursting_master_requests = cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;

  //clock_crossing_ddr2_cpu_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_any_bursting_master_saved_grant = 0;

  //clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value = clock_crossing_ddr2_cpu_s1_firsttransfer ? (clock_crossing_ddr2_cpu_s1_arb_share_set_values - 1) : |clock_crossing_ddr2_cpu_s1_arb_share_counter ? (clock_crossing_ddr2_cpu_s1_arb_share_counter - 1) : 0;

  //clock_crossing_ddr2_cpu_s1_allgrants all slave grants, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_allgrants = |clock_crossing_ddr2_cpu_s1_grant_vector;

  //clock_crossing_ddr2_cpu_s1_end_xfer assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_end_xfer = ~(clock_crossing_ddr2_cpu_s1_waits_for_read | clock_crossing_ddr2_cpu_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1 = clock_crossing_ddr2_cpu_s1_end_xfer & (~clock_crossing_ddr2_cpu_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //clock_crossing_ddr2_cpu_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1 & clock_crossing_ddr2_cpu_s1_allgrants) | (end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1 & ~clock_crossing_ddr2_cpu_s1_non_bursting_master_requests);

  //clock_crossing_ddr2_cpu_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_s1_arb_share_counter <= 0;
      else if (clock_crossing_ddr2_cpu_s1_arb_counter_enable)
          clock_crossing_ddr2_cpu_s1_arb_share_counter <= clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value;
    end


  //clock_crossing_ddr2_cpu_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_s1_slavearbiterlockenable <= 0;
      else if ((|clock_crossing_ddr2_cpu_s1_master_qreq_vector & end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1) | (end_xfer_arb_share_counter_term_clock_crossing_ddr2_cpu_s1 & ~clock_crossing_ddr2_cpu_s1_non_bursting_master_requests))
          clock_crossing_ddr2_cpu_s1_slavearbiterlockenable <= |clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value;
    end


  //cpu/data_master clock_crossing_ddr2_cpu/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = clock_crossing_ddr2_cpu_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //clock_crossing_ddr2_cpu_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_slavearbiterlockenable2 = |clock_crossing_ddr2_cpu_s1_arb_share_counter_next_value;

  //cpu/data_master clock_crossing_ddr2_cpu/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = clock_crossing_ddr2_cpu_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //clock_crossing_ddr2_cpu_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1 = cpu_data_master_requests_clock_crossing_ddr2_cpu_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter))));
  //unique name for clock_crossing_ddr2_cpu_s1_move_on_to_next_transaction, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_move_on_to_next_transaction = clock_crossing_ddr2_cpu_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_clock_crossing_ddr2_cpu_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_clock_crossing_ddr2_cpu_s1_module rdv_fifo_for_cpu_data_master_to_clock_crossing_ddr2_cpu_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_clock_crossing_ddr2_cpu_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_clock_crossing_ddr2_cpu_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_clock_crossing_ddr2_cpu_s1),
      .full                 (),
      .read                 (clock_crossing_ddr2_cpu_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_ddr2_cpu_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_clock_crossing_ddr2_cpu_s1;
  //local readdatavalid cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1 = clock_crossing_ddr2_cpu_s1_readdatavalid_from_sa;

  //clock_crossing_ddr2_cpu_s1_writedata mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_writedata = cpu_data_master_writedata;

  //assign clock_crossing_ddr2_cpu_s1_endofpacket_from_sa = clock_crossing_ddr2_cpu_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_endofpacket_from_sa = clock_crossing_ddr2_cpu_s1_endofpacket;

  //master is always granted when requested
  assign cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 = cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1;

  //cpu/data_master saved-grant clock_crossing_ddr2_cpu/s1, which is an e_assign
  assign cpu_data_master_saved_grant_clock_crossing_ddr2_cpu_s1 = cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;

  //allow new arb cycle for clock_crossing_ddr2_cpu/s1, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign clock_crossing_ddr2_cpu_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign clock_crossing_ddr2_cpu_s1_master_qreq_vector = 1;

  //clock_crossing_ddr2_cpu_s1_reset_n assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_reset_n = reset_n;

  //clock_crossing_ddr2_cpu_s1_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_firsttransfer = clock_crossing_ddr2_cpu_s1_begins_xfer ? clock_crossing_ddr2_cpu_s1_unreg_firsttransfer : clock_crossing_ddr2_cpu_s1_reg_firsttransfer;

  //clock_crossing_ddr2_cpu_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_unreg_firsttransfer = ~(clock_crossing_ddr2_cpu_s1_slavearbiterlockenable & clock_crossing_ddr2_cpu_s1_any_continuerequest);

  //clock_crossing_ddr2_cpu_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_s1_reg_firsttransfer <= 1'b1;
      else if (clock_crossing_ddr2_cpu_s1_begins_xfer)
          clock_crossing_ddr2_cpu_s1_reg_firsttransfer <= clock_crossing_ddr2_cpu_s1_unreg_firsttransfer;
    end


  //clock_crossing_ddr2_cpu_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_beginbursttransfer_internal = clock_crossing_ddr2_cpu_s1_begins_xfer;

  //clock_crossing_ddr2_cpu_s1_read assignment, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_read = cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 & cpu_data_master_read;

  //clock_crossing_ddr2_cpu_s1_write assignment, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_write = cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 & cpu_data_master_write;

  assign shifted_address_to_clock_crossing_ddr2_cpu_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //clock_crossing_ddr2_cpu_s1_address mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_address = shifted_address_to_clock_crossing_ddr2_cpu_s1_from_cpu_data_master >> 2;

  //slaveid clock_crossing_ddr2_cpu_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_nativeaddress = cpu_data_master_address_to_slave >> 2;

  //d1_clock_crossing_ddr2_cpu_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_clock_crossing_ddr2_cpu_s1_end_xfer <= 1;
      else 
        d1_clock_crossing_ddr2_cpu_s1_end_xfer <= clock_crossing_ddr2_cpu_s1_end_xfer;
    end


  //clock_crossing_ddr2_cpu_s1_waits_for_read in a cycle, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_waits_for_read = clock_crossing_ddr2_cpu_s1_in_a_read_cycle & clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;

  //clock_crossing_ddr2_cpu_s1_in_a_read_cycle assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_in_a_read_cycle = cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = clock_crossing_ddr2_cpu_s1_in_a_read_cycle;

  //clock_crossing_ddr2_cpu_s1_waits_for_write in a cycle, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_waits_for_write = clock_crossing_ddr2_cpu_s1_in_a_write_cycle & clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;

  //clock_crossing_ddr2_cpu_s1_in_a_write_cycle assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_s1_in_a_write_cycle = cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = clock_crossing_ddr2_cpu_s1_in_a_write_cycle;

  assign wait_for_clock_crossing_ddr2_cpu_s1_counter = 0;
  //clock_crossing_ddr2_cpu_s1_byteenable byte enable port mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_s1_byteenable = (cpu_data_master_granted_clock_crossing_ddr2_cpu_s1)? cpu_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_ddr2_cpu/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_ddr2_cpu_m1_arbitrator (
                                               // inputs:
                                                clk,
                                                clock_crossing_ddr2_cpu_m1_address,
                                                clock_crossing_ddr2_cpu_m1_byteenable,
                                                clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1,
                                                clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1,
                                                clock_crossing_ddr2_cpu_m1_read,
                                                clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1,
                                                clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register,
                                                clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1,
                                                clock_crossing_ddr2_cpu_m1_write,
                                                clock_crossing_ddr2_cpu_m1_writedata,
                                                d1_pipeline_bridge_ddr2_s1_end_xfer,
                                                pipeline_bridge_ddr2_s1_endofpacket_from_sa,
                                                pipeline_bridge_ddr2_s1_readdata_from_sa,
                                                pipeline_bridge_ddr2_s1_waitrequest_from_sa,
                                                reset_n,

                                               // outputs:
                                                clock_crossing_ddr2_cpu_m1_address_to_slave,
                                                clock_crossing_ddr2_cpu_m1_endofpacket,
                                                clock_crossing_ddr2_cpu_m1_latency_counter,
                                                clock_crossing_ddr2_cpu_m1_readdata,
                                                clock_crossing_ddr2_cpu_m1_readdatavalid,
                                                clock_crossing_ddr2_cpu_m1_reset_n,
                                                clock_crossing_ddr2_cpu_m1_waitrequest
                                             )
;

  output  [ 29: 0] clock_crossing_ddr2_cpu_m1_address_to_slave;
  output           clock_crossing_ddr2_cpu_m1_endofpacket;
  output           clock_crossing_ddr2_cpu_m1_latency_counter;
  output  [ 31: 0] clock_crossing_ddr2_cpu_m1_readdata;
  output           clock_crossing_ddr2_cpu_m1_readdatavalid;
  output           clock_crossing_ddr2_cpu_m1_reset_n;
  output           clock_crossing_ddr2_cpu_m1_waitrequest;
  input            clk;
  input   [ 29: 0] clock_crossing_ddr2_cpu_m1_address;
  input   [  3: 0] clock_crossing_ddr2_cpu_m1_byteenable;
  input            clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1;
  input            clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1;
  input            clock_crossing_ddr2_cpu_m1_read;
  input            clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1;
  input            clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register;
  input            clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;
  input            clock_crossing_ddr2_cpu_m1_write;
  input   [ 31: 0] clock_crossing_ddr2_cpu_m1_writedata;
  input            d1_pipeline_bridge_ddr2_s1_end_xfer;
  input            pipeline_bridge_ddr2_s1_endofpacket_from_sa;
  input   [ 31: 0] pipeline_bridge_ddr2_s1_readdata_from_sa;
  input            pipeline_bridge_ddr2_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 29: 0] clock_crossing_ddr2_cpu_m1_address_last_time;
  wire    [ 29: 0] clock_crossing_ddr2_cpu_m1_address_to_slave;
  reg     [  3: 0] clock_crossing_ddr2_cpu_m1_byteenable_last_time;
  wire             clock_crossing_ddr2_cpu_m1_endofpacket;
  wire             clock_crossing_ddr2_cpu_m1_latency_counter;
  reg              clock_crossing_ddr2_cpu_m1_read_last_time;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_m1_readdata;
  wire             clock_crossing_ddr2_cpu_m1_readdatavalid;
  wire             clock_crossing_ddr2_cpu_m1_reset_n;
  wire             clock_crossing_ddr2_cpu_m1_run;
  wire             clock_crossing_ddr2_cpu_m1_waitrequest;
  reg              clock_crossing_ddr2_cpu_m1_write_last_time;
  reg     [ 31: 0] clock_crossing_ddr2_cpu_m1_writedata_last_time;
  wire             pre_flush_clock_crossing_ddr2_cpu_m1_readdatavalid;
  wire             r_2;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1 | ~clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1) & ((~clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1 | ~(clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write) | (1 & ~pipeline_bridge_ddr2_s1_waitrequest_from_sa & (clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write)))) & ((~clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1 | ~(clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write) | (1 & ~pipeline_bridge_ddr2_s1_waitrequest_from_sa & (clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write))));

  //cascaded wait assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign clock_crossing_ddr2_cpu_m1_address_to_slave = clock_crossing_ddr2_cpu_m1_address[29 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_clock_crossing_ddr2_cpu_m1_readdatavalid = clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign clock_crossing_ddr2_cpu_m1_readdatavalid = 0 |
    pre_flush_clock_crossing_ddr2_cpu_m1_readdatavalid;

  //clock_crossing_ddr2_cpu/m1 readdata mux, which is an e_mux
  assign clock_crossing_ddr2_cpu_m1_readdata = pipeline_bridge_ddr2_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_waitrequest = ~clock_crossing_ddr2_cpu_m1_run;

  //latent max counter, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_latency_counter = 0;

  //clock_crossing_ddr2_cpu_m1_reset_n assignment, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_reset_n = reset_n;

  //mux clock_crossing_ddr2_cpu_m1_endofpacket, which is an e_mux
  assign clock_crossing_ddr2_cpu_m1_endofpacket = pipeline_bridge_ddr2_s1_endofpacket_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_ddr2_cpu_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_m1_address_last_time <= 0;
      else 
        clock_crossing_ddr2_cpu_m1_address_last_time <= clock_crossing_ddr2_cpu_m1_address;
    end


  //clock_crossing_ddr2_cpu/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= clock_crossing_ddr2_cpu_m1_waitrequest & (clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write);
    end


  //clock_crossing_ddr2_cpu_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_ddr2_cpu_m1_address != clock_crossing_ddr2_cpu_m1_address_last_time))
        begin
          $write("%0d ns: clock_crossing_ddr2_cpu_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_ddr2_cpu_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_m1_byteenable_last_time <= 0;
      else 
        clock_crossing_ddr2_cpu_m1_byteenable_last_time <= clock_crossing_ddr2_cpu_m1_byteenable;
    end


  //clock_crossing_ddr2_cpu_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_ddr2_cpu_m1_byteenable != clock_crossing_ddr2_cpu_m1_byteenable_last_time))
        begin
          $write("%0d ns: clock_crossing_ddr2_cpu_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_ddr2_cpu_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_m1_read_last_time <= 0;
      else 
        clock_crossing_ddr2_cpu_m1_read_last_time <= clock_crossing_ddr2_cpu_m1_read;
    end


  //clock_crossing_ddr2_cpu_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_ddr2_cpu_m1_read != clock_crossing_ddr2_cpu_m1_read_last_time))
        begin
          $write("%0d ns: clock_crossing_ddr2_cpu_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_ddr2_cpu_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_m1_write_last_time <= 0;
      else 
        clock_crossing_ddr2_cpu_m1_write_last_time <= clock_crossing_ddr2_cpu_m1_write;
    end


  //clock_crossing_ddr2_cpu_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_ddr2_cpu_m1_write != clock_crossing_ddr2_cpu_m1_write_last_time))
        begin
          $write("%0d ns: clock_crossing_ddr2_cpu_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_ddr2_cpu_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_ddr2_cpu_m1_writedata_last_time <= 0;
      else 
        clock_crossing_ddr2_cpu_m1_writedata_last_time <= clock_crossing_ddr2_cpu_m1_writedata;
    end


  //clock_crossing_ddr2_cpu_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_ddr2_cpu_m1_writedata != clock_crossing_ddr2_cpu_m1_writedata_last_time) & clock_crossing_ddr2_cpu_m1_write)
        begin
          $write("%0d ns: clock_crossing_ddr2_cpu_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_ddr2_cpu_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_clock_crossing_master_ddr2_s1_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  3: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  3: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  3: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  3: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  3: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  3: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  3: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  3: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  3: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  3: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  3: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  3: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  3: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  3: 0] p31_stage_31;
  wire             p32_full_32;
  wire    [  3: 0] p32_stage_32;
  wire             p33_full_33;
  wire    [  3: 0] p33_stage_33;
  wire             p34_full_34;
  wire    [  3: 0] p34_stage_34;
  wire             p35_full_35;
  wire    [  3: 0] p35_stage_35;
  wire             p36_full_36;
  wire    [  3: 0] p36_stage_36;
  wire             p37_full_37;
  wire    [  3: 0] p37_stage_37;
  wire             p38_full_38;
  wire    [  3: 0] p38_stage_38;
  wire             p39_full_39;
  wire    [  3: 0] p39_stage_39;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p40_full_40;
  wire    [  3: 0] p40_stage_40;
  wire             p41_full_41;
  wire    [  3: 0] p41_stage_41;
  wire             p42_full_42;
  wire    [  3: 0] p42_stage_42;
  wire             p43_full_43;
  wire    [  3: 0] p43_stage_43;
  wire             p44_full_44;
  wire    [  3: 0] p44_stage_44;
  wire             p45_full_45;
  wire    [  3: 0] p45_stage_45;
  wire             p46_full_46;
  wire    [  3: 0] p46_stage_46;
  wire             p47_full_47;
  wire    [  3: 0] p47_stage_47;
  wire             p48_full_48;
  wire    [  3: 0] p48_stage_48;
  wire             p49_full_49;
  wire    [  3: 0] p49_stage_49;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p50_full_50;
  wire    [  3: 0] p50_stage_50;
  wire             p51_full_51;
  wire    [  3: 0] p51_stage_51;
  wire             p52_full_52;
  wire    [  3: 0] p52_stage_52;
  wire             p53_full_53;
  wire    [  3: 0] p53_stage_53;
  wire             p54_full_54;
  wire    [  3: 0] p54_stage_54;
  wire             p55_full_55;
  wire    [  3: 0] p55_stage_55;
  wire             p56_full_56;
  wire    [  3: 0] p56_stage_56;
  wire             p57_full_57;
  wire    [  3: 0] p57_stage_57;
  wire             p58_full_58;
  wire    [  3: 0] p58_stage_58;
  wire             p59_full_59;
  wire    [  3: 0] p59_stage_59;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p60_full_60;
  wire    [  3: 0] p60_stage_60;
  wire             p61_full_61;
  wire    [  3: 0] p61_stage_61;
  wire             p62_full_62;
  wire    [  3: 0] p62_stage_62;
  wire             p63_full_63;
  wire    [  3: 0] p63_stage_63;
  wire             p64_full_64;
  wire    [  3: 0] p64_stage_64;
  wire             p65_full_65;
  wire    [  3: 0] p65_stage_65;
  wire             p66_full_66;
  wire    [  3: 0] p66_stage_66;
  wire             p67_full_67;
  wire    [  3: 0] p67_stage_67;
  wire             p68_full_68;
  wire    [  3: 0] p68_stage_68;
  wire             p69_full_69;
  wire    [  3: 0] p69_stage_69;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p70_full_70;
  wire    [  3: 0] p70_stage_70;
  wire             p71_full_71;
  wire    [  3: 0] p71_stage_71;
  wire             p72_full_72;
  wire    [  3: 0] p72_stage_72;
  wire             p73_full_73;
  wire    [  3: 0] p73_stage_73;
  wire             p74_full_74;
  wire    [  3: 0] p74_stage_74;
  wire             p75_full_75;
  wire    [  3: 0] p75_stage_75;
  wire             p76_full_76;
  wire    [  3: 0] p76_stage_76;
  wire             p77_full_77;
  wire    [  3: 0] p77_stage_77;
  wire             p78_full_78;
  wire    [  3: 0] p78_stage_78;
  wire             p79_full_79;
  wire    [  3: 0] p79_stage_79;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p80_full_80;
  wire    [  3: 0] p80_stage_80;
  wire             p81_full_81;
  wire    [  3: 0] p81_stage_81;
  wire             p82_full_82;
  wire    [  3: 0] p82_stage_82;
  wire             p83_full_83;
  wire    [  3: 0] p83_stage_83;
  wire             p84_full_84;
  wire    [  3: 0] p84_stage_84;
  wire             p85_full_85;
  wire    [  3: 0] p85_stage_85;
  wire             p86_full_86;
  wire    [  3: 0] p86_stage_86;
  wire             p87_full_87;
  wire    [  3: 0] p87_stage_87;
  wire             p88_full_88;
  wire    [  3: 0] p88_stage_88;
  wire             p89_full_89;
  wire    [  3: 0] p89_stage_89;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p90_full_90;
  wire    [  3: 0] p90_stage_90;
  wire             p91_full_91;
  wire    [  3: 0] p91_stage_91;
  wire             p92_full_92;
  wire    [  3: 0] p92_stage_92;
  wire             p93_full_93;
  wire    [  3: 0] p93_stage_93;
  wire             p94_full_94;
  wire    [  3: 0] p94_stage_94;
  wire             p95_full_95;
  wire    [  3: 0] p95_stage_95;
  wire             p96_full_96;
  wire    [  3: 0] p96_stage_96;
  wire             p97_full_97;
  wire    [  3: 0] p97_stage_97;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_18;
  reg     [  3: 0] stage_19;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_20;
  reg     [  3: 0] stage_21;
  reg     [  3: 0] stage_22;
  reg     [  3: 0] stage_23;
  reg     [  3: 0] stage_24;
  reg     [  3: 0] stage_25;
  reg     [  3: 0] stage_26;
  reg     [  3: 0] stage_27;
  reg     [  3: 0] stage_28;
  reg     [  3: 0] stage_29;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_30;
  reg     [  3: 0] stage_31;
  reg     [  3: 0] stage_32;
  reg     [  3: 0] stage_33;
  reg     [  3: 0] stage_34;
  reg     [  3: 0] stage_35;
  reg     [  3: 0] stage_36;
  reg     [  3: 0] stage_37;
  reg     [  3: 0] stage_38;
  reg     [  3: 0] stage_39;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_40;
  reg     [  3: 0] stage_41;
  reg     [  3: 0] stage_42;
  reg     [  3: 0] stage_43;
  reg     [  3: 0] stage_44;
  reg     [  3: 0] stage_45;
  reg     [  3: 0] stage_46;
  reg     [  3: 0] stage_47;
  reg     [  3: 0] stage_48;
  reg     [  3: 0] stage_49;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_50;
  reg     [  3: 0] stage_51;
  reg     [  3: 0] stage_52;
  reg     [  3: 0] stage_53;
  reg     [  3: 0] stage_54;
  reg     [  3: 0] stage_55;
  reg     [  3: 0] stage_56;
  reg     [  3: 0] stage_57;
  reg     [  3: 0] stage_58;
  reg     [  3: 0] stage_59;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_60;
  reg     [  3: 0] stage_61;
  reg     [  3: 0] stage_62;
  reg     [  3: 0] stage_63;
  reg     [  3: 0] stage_64;
  reg     [  3: 0] stage_65;
  reg     [  3: 0] stage_66;
  reg     [  3: 0] stage_67;
  reg     [  3: 0] stage_68;
  reg     [  3: 0] stage_69;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_70;
  reg     [  3: 0] stage_71;
  reg     [  3: 0] stage_72;
  reg     [  3: 0] stage_73;
  reg     [  3: 0] stage_74;
  reg     [  3: 0] stage_75;
  reg     [  3: 0] stage_76;
  reg     [  3: 0] stage_77;
  reg     [  3: 0] stage_78;
  reg     [  3: 0] stage_79;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_80;
  reg     [  3: 0] stage_81;
  reg     [  3: 0] stage_82;
  reg     [  3: 0] stage_83;
  reg     [  3: 0] stage_84;
  reg     [  3: 0] stage_85;
  reg     [  3: 0] stage_86;
  reg     [  3: 0] stage_87;
  reg     [  3: 0] stage_88;
  reg     [  3: 0] stage_89;
  reg     [  3: 0] stage_9;
  reg     [  3: 0] stage_90;
  reg     [  3: 0] stage_91;
  reg     [  3: 0] stage_92;
  reg     [  3: 0] stage_93;
  reg     [  3: 0] stage_94;
  reg     [  3: 0] stage_95;
  reg     [  3: 0] stage_96;
  reg     [  3: 0] stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_master_read_avalon_master_to_clock_crossing_master_ddr2_s1_module (
                                                                                        // inputs:
                                                                                         clear_fifo,
                                                                                         clk,
                                                                                         data_in,
                                                                                         read,
                                                                                         reset_n,
                                                                                         sync_reset,
                                                                                         write,

                                                                                        // outputs:
                                                                                         data_out,
                                                                                         empty,
                                                                                         fifo_contains_ones_n,
                                                                                         full
                                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p96_full_96;
  wire             p96_stage_96;
  wire             p97_full_97;
  wire             p97_stage_97;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  reg              stage_96;
  reg              stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_master_ddr2_s1_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   clock_crossing_master_ddr2_s1_endofpacket,
                                                   clock_crossing_master_ddr2_s1_readdata,
                                                   clock_crossing_master_ddr2_s1_readdatavalid,
                                                   clock_crossing_master_ddr2_s1_waitrequest,
                                                   master_read_avalon_master_address_to_slave,
                                                   master_read_avalon_master_burstcount,
                                                   master_read_avalon_master_read,
                                                   master_read_latency_counter,
                                                   master_write_avalon_master_address_to_slave,
                                                   master_write_avalon_master_burstcount,
                                                   master_write_avalon_master_byteenable,
                                                   master_write_avalon_master_write,
                                                   master_write_avalon_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   clock_crossing_master_ddr2_s1_address,
                                                   clock_crossing_master_ddr2_s1_burstcount,
                                                   clock_crossing_master_ddr2_s1_byteenable,
                                                   clock_crossing_master_ddr2_s1_endofpacket_from_sa,
                                                   clock_crossing_master_ddr2_s1_nativeaddress,
                                                   clock_crossing_master_ddr2_s1_read,
                                                   clock_crossing_master_ddr2_s1_readdata_from_sa,
                                                   clock_crossing_master_ddr2_s1_reset_n,
                                                   clock_crossing_master_ddr2_s1_waitrequest_from_sa,
                                                   clock_crossing_master_ddr2_s1_write,
                                                   clock_crossing_master_ddr2_s1_writedata,
                                                   d1_clock_crossing_master_ddr2_s1_end_xfer,
                                                   master_read_granted_clock_crossing_master_ddr2_s1,
                                                   master_read_qualified_request_clock_crossing_master_ddr2_s1,
                                                   master_read_read_data_valid_clock_crossing_master_ddr2_s1,
                                                   master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register,
                                                   master_read_requests_clock_crossing_master_ddr2_s1,
                                                   master_write_granted_clock_crossing_master_ddr2_s1,
                                                   master_write_qualified_request_clock_crossing_master_ddr2_s1,
                                                   master_write_requests_clock_crossing_master_ddr2_s1
                                                )
;

  output  [ 24: 0] clock_crossing_master_ddr2_s1_address;
  output  [  3: 0] clock_crossing_master_ddr2_s1_burstcount;
  output  [ 31: 0] clock_crossing_master_ddr2_s1_byteenable;
  output           clock_crossing_master_ddr2_s1_endofpacket_from_sa;
  output  [ 24: 0] clock_crossing_master_ddr2_s1_nativeaddress;
  output           clock_crossing_master_ddr2_s1_read;
  output  [255: 0] clock_crossing_master_ddr2_s1_readdata_from_sa;
  output           clock_crossing_master_ddr2_s1_reset_n;
  output           clock_crossing_master_ddr2_s1_waitrequest_from_sa;
  output           clock_crossing_master_ddr2_s1_write;
  output  [255: 0] clock_crossing_master_ddr2_s1_writedata;
  output           d1_clock_crossing_master_ddr2_s1_end_xfer;
  output           master_read_granted_clock_crossing_master_ddr2_s1;
  output           master_read_qualified_request_clock_crossing_master_ddr2_s1;
  output           master_read_read_data_valid_clock_crossing_master_ddr2_s1;
  output           master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register;
  output           master_read_requests_clock_crossing_master_ddr2_s1;
  output           master_write_granted_clock_crossing_master_ddr2_s1;
  output           master_write_qualified_request_clock_crossing_master_ddr2_s1;
  output           master_write_requests_clock_crossing_master_ddr2_s1;
  input            clk;
  input            clock_crossing_master_ddr2_s1_endofpacket;
  input   [255: 0] clock_crossing_master_ddr2_s1_readdata;
  input            clock_crossing_master_ddr2_s1_readdatavalid;
  input            clock_crossing_master_ddr2_s1_waitrequest;
  input   [ 29: 0] master_read_avalon_master_address_to_slave;
  input   [  3: 0] master_read_avalon_master_burstcount;
  input            master_read_avalon_master_read;
  input            master_read_latency_counter;
  input   [ 29: 0] master_write_avalon_master_address_to_slave;
  input   [  3: 0] master_write_avalon_master_burstcount;
  input   [ 31: 0] master_write_avalon_master_byteenable;
  input            master_write_avalon_master_write;
  input   [255: 0] master_write_avalon_master_writedata;
  input            reset_n;

  wire    [ 24: 0] clock_crossing_master_ddr2_s1_address;
  wire             clock_crossing_master_ddr2_s1_allgrants;
  wire             clock_crossing_master_ddr2_s1_allow_new_arb_cycle;
  wire             clock_crossing_master_ddr2_s1_any_bursting_master_saved_grant;
  wire             clock_crossing_master_ddr2_s1_any_continuerequest;
  reg     [  1: 0] clock_crossing_master_ddr2_s1_arb_addend;
  wire             clock_crossing_master_ddr2_s1_arb_counter_enable;
  reg     [  3: 0] clock_crossing_master_ddr2_s1_arb_share_counter;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_arb_share_counter_next_value;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_arb_share_set_values;
  wire    [  1: 0] clock_crossing_master_ddr2_s1_arb_winner;
  wire             clock_crossing_master_ddr2_s1_arbitration_holdoff_internal;
  reg     [  2: 0] clock_crossing_master_ddr2_s1_bbt_burstcounter;
  wire             clock_crossing_master_ddr2_s1_beginbursttransfer_internal;
  wire             clock_crossing_master_ddr2_s1_begins_xfer;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_burstcount;
  wire             clock_crossing_master_ddr2_s1_burstcount_fifo_empty;
  wire    [ 31: 0] clock_crossing_master_ddr2_s1_byteenable;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_chosen_master_double_vector;
  wire    [  1: 0] clock_crossing_master_ddr2_s1_chosen_master_rot_left;
  reg     [  3: 0] clock_crossing_master_ddr2_s1_current_burst;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_current_burst_minus_one;
  wire             clock_crossing_master_ddr2_s1_end_xfer;
  wire             clock_crossing_master_ddr2_s1_endofpacket_from_sa;
  wire             clock_crossing_master_ddr2_s1_firsttransfer;
  wire    [  1: 0] clock_crossing_master_ddr2_s1_grant_vector;
  wire             clock_crossing_master_ddr2_s1_in_a_read_cycle;
  wire             clock_crossing_master_ddr2_s1_in_a_write_cycle;
  reg              clock_crossing_master_ddr2_s1_load_fifo;
  wire    [  1: 0] clock_crossing_master_ddr2_s1_master_qreq_vector;
  wire             clock_crossing_master_ddr2_s1_move_on_to_next_transaction;
  wire    [ 24: 0] clock_crossing_master_ddr2_s1_nativeaddress;
  wire    [  2: 0] clock_crossing_master_ddr2_s1_next_bbt_burstcount;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_next_burst_count;
  wire             clock_crossing_master_ddr2_s1_non_bursting_master_requests;
  wire             clock_crossing_master_ddr2_s1_read;
  wire    [255: 0] clock_crossing_master_ddr2_s1_readdata_from_sa;
  wire             clock_crossing_master_ddr2_s1_readdatavalid_from_sa;
  reg              clock_crossing_master_ddr2_s1_reg_firsttransfer;
  wire             clock_crossing_master_ddr2_s1_reset_n;
  reg     [  1: 0] clock_crossing_master_ddr2_s1_saved_chosen_master_vector;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_selected_burstcount;
  reg              clock_crossing_master_ddr2_s1_slavearbiterlockenable;
  wire             clock_crossing_master_ddr2_s1_slavearbiterlockenable2;
  wire             clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_transaction_burst_count;
  wire             clock_crossing_master_ddr2_s1_unreg_firsttransfer;
  wire             clock_crossing_master_ddr2_s1_waitrequest_from_sa;
  wire             clock_crossing_master_ddr2_s1_waits_for_read;
  wire             clock_crossing_master_ddr2_s1_waits_for_write;
  wire             clock_crossing_master_ddr2_s1_write;
  wire    [255: 0] clock_crossing_master_ddr2_s1_writedata;
  reg              d1_clock_crossing_master_ddr2_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_master_read_avalon_master_granted_slave_clock_crossing_master_ddr2_s1;
  reg              last_cycle_master_write_avalon_master_granted_slave_clock_crossing_master_ddr2_s1;
  wire             master_read_avalon_master_arbiterlock;
  wire             master_read_avalon_master_arbiterlock2;
  wire             master_read_avalon_master_continuerequest;
  wire             master_read_granted_clock_crossing_master_ddr2_s1;
  wire             master_read_qualified_request_clock_crossing_master_ddr2_s1;
  wire             master_read_rdv_fifo_empty_clock_crossing_master_ddr2_s1;
  wire             master_read_rdv_fifo_output_from_clock_crossing_master_ddr2_s1;
  wire             master_read_read_data_valid_clock_crossing_master_ddr2_s1;
  wire             master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register;
  wire             master_read_requests_clock_crossing_master_ddr2_s1;
  wire             master_read_saved_grant_clock_crossing_master_ddr2_s1;
  wire             master_write_avalon_master_arbiterlock;
  wire             master_write_avalon_master_arbiterlock2;
  wire             master_write_avalon_master_continuerequest;
  wire             master_write_granted_clock_crossing_master_ddr2_s1;
  wire             master_write_qualified_request_clock_crossing_master_ddr2_s1;
  wire             master_write_requests_clock_crossing_master_ddr2_s1;
  wire             master_write_saved_grant_clock_crossing_master_ddr2_s1;
  wire             p0_clock_crossing_master_ddr2_s1_load_fifo;
  wire    [ 29: 0] shifted_address_to_clock_crossing_master_ddr2_s1_from_master_read_avalon_master;
  wire    [ 29: 0] shifted_address_to_clock_crossing_master_ddr2_s1_from_master_write_avalon_master;
  wire             wait_for_clock_crossing_master_ddr2_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~clock_crossing_master_ddr2_s1_end_xfer;
    end


  assign clock_crossing_master_ddr2_s1_begins_xfer = ~d1_reasons_to_wait & ((master_read_qualified_request_clock_crossing_master_ddr2_s1 | master_write_qualified_request_clock_crossing_master_ddr2_s1));
  //assign clock_crossing_master_ddr2_s1_readdata_from_sa = clock_crossing_master_ddr2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_master_ddr2_s1_readdata_from_sa = clock_crossing_master_ddr2_s1_readdata;

  assign master_read_requests_clock_crossing_master_ddr2_s1 = ((1) & (master_read_avalon_master_read)) & master_read_avalon_master_read;
  //assign clock_crossing_master_ddr2_s1_waitrequest_from_sa = clock_crossing_master_ddr2_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_master_ddr2_s1_waitrequest_from_sa = clock_crossing_master_ddr2_s1_waitrequest;

  //assign clock_crossing_master_ddr2_s1_readdatavalid_from_sa = clock_crossing_master_ddr2_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_master_ddr2_s1_readdatavalid_from_sa = clock_crossing_master_ddr2_s1_readdatavalid;

  //clock_crossing_master_ddr2_s1_arb_share_counter set values, which is an e_mux
  assign clock_crossing_master_ddr2_s1_arb_share_set_values = (master_write_granted_clock_crossing_master_ddr2_s1)? master_write_avalon_master_burstcount :
    (master_write_granted_clock_crossing_master_ddr2_s1)? master_write_avalon_master_burstcount :
    1;

  //clock_crossing_master_ddr2_s1_non_bursting_master_requests mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_non_bursting_master_requests = 0;

  //clock_crossing_master_ddr2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_any_bursting_master_saved_grant = master_read_saved_grant_clock_crossing_master_ddr2_s1 |
    master_write_saved_grant_clock_crossing_master_ddr2_s1 |
    master_read_saved_grant_clock_crossing_master_ddr2_s1 |
    master_write_saved_grant_clock_crossing_master_ddr2_s1;

  //clock_crossing_master_ddr2_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign clock_crossing_master_ddr2_s1_arb_share_counter_next_value = clock_crossing_master_ddr2_s1_firsttransfer ? (clock_crossing_master_ddr2_s1_arb_share_set_values - 1) : |clock_crossing_master_ddr2_s1_arb_share_counter ? (clock_crossing_master_ddr2_s1_arb_share_counter - 1) : 0;

  //clock_crossing_master_ddr2_s1_allgrants all slave grants, which is an e_mux
  assign clock_crossing_master_ddr2_s1_allgrants = (|clock_crossing_master_ddr2_s1_grant_vector) |
    (|clock_crossing_master_ddr2_s1_grant_vector) |
    (|clock_crossing_master_ddr2_s1_grant_vector) |
    (|clock_crossing_master_ddr2_s1_grant_vector);

  //clock_crossing_master_ddr2_s1_end_xfer assignment, which is an e_assign
  assign clock_crossing_master_ddr2_s1_end_xfer = ~(clock_crossing_master_ddr2_s1_waits_for_read | clock_crossing_master_ddr2_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1 = clock_crossing_master_ddr2_s1_end_xfer & (~clock_crossing_master_ddr2_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //clock_crossing_master_ddr2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign clock_crossing_master_ddr2_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1 & clock_crossing_master_ddr2_s1_allgrants) | (end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1 & ~clock_crossing_master_ddr2_s1_non_bursting_master_requests);

  //clock_crossing_master_ddr2_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_arb_share_counter <= 0;
      else if (clock_crossing_master_ddr2_s1_arb_counter_enable)
          clock_crossing_master_ddr2_s1_arb_share_counter <= clock_crossing_master_ddr2_s1_arb_share_counter_next_value;
    end


  //clock_crossing_master_ddr2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_slavearbiterlockenable <= 0;
      else if ((|clock_crossing_master_ddr2_s1_master_qreq_vector & end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1) | (end_xfer_arb_share_counter_term_clock_crossing_master_ddr2_s1 & ~clock_crossing_master_ddr2_s1_non_bursting_master_requests))
          clock_crossing_master_ddr2_s1_slavearbiterlockenable <= |clock_crossing_master_ddr2_s1_arb_share_counter_next_value;
    end


  //master_read/avalon_master clock_crossing_master_ddr2/s1 arbiterlock, which is an e_assign
  assign master_read_avalon_master_arbiterlock = clock_crossing_master_ddr2_s1_slavearbiterlockenable & master_read_avalon_master_continuerequest;

  //clock_crossing_master_ddr2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign clock_crossing_master_ddr2_s1_slavearbiterlockenable2 = |clock_crossing_master_ddr2_s1_arb_share_counter_next_value;

  //master_read/avalon_master clock_crossing_master_ddr2/s1 arbiterlock2, which is an e_assign
  assign master_read_avalon_master_arbiterlock2 = clock_crossing_master_ddr2_s1_slavearbiterlockenable2 & master_read_avalon_master_continuerequest;

  //master_write/avalon_master clock_crossing_master_ddr2/s1 arbiterlock, which is an e_assign
  assign master_write_avalon_master_arbiterlock = clock_crossing_master_ddr2_s1_slavearbiterlockenable & master_write_avalon_master_continuerequest;

  //master_write/avalon_master clock_crossing_master_ddr2/s1 arbiterlock2, which is an e_assign
  assign master_write_avalon_master_arbiterlock2 = clock_crossing_master_ddr2_s1_slavearbiterlockenable2 & master_write_avalon_master_continuerequest;

  //master_write/avalon_master granted clock_crossing_master_ddr2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_master_write_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 <= 0;
      else 
        last_cycle_master_write_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 <= master_write_saved_grant_clock_crossing_master_ddr2_s1 ? 1 : (clock_crossing_master_ddr2_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_master_write_avalon_master_granted_slave_clock_crossing_master_ddr2_s1;
    end


  //master_write_avalon_master_continuerequest continued request, which is an e_mux
  assign master_write_avalon_master_continuerequest = last_cycle_master_write_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 & 1;

  //clock_crossing_master_ddr2_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign clock_crossing_master_ddr2_s1_any_continuerequest = master_write_avalon_master_continuerequest |
    master_read_avalon_master_continuerequest;

  assign master_read_qualified_request_clock_crossing_master_ddr2_s1 = master_read_requests_clock_crossing_master_ddr2_s1 & ~((master_read_avalon_master_read & ((master_read_latency_counter != 0) | (1 < master_read_latency_counter))) | master_write_avalon_master_arbiterlock);
  //unique name for clock_crossing_master_ddr2_s1_move_on_to_next_transaction, which is an e_assign
  assign clock_crossing_master_ddr2_s1_move_on_to_next_transaction = clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst & clock_crossing_master_ddr2_s1_load_fifo;

  //the currently selected burstcount for clock_crossing_master_ddr2_s1, which is an e_mux
  assign clock_crossing_master_ddr2_s1_selected_burstcount = (master_read_granted_clock_crossing_master_ddr2_s1)? master_read_avalon_master_burstcount :
    1;

  //burstcount_fifo_for_clock_crossing_master_ddr2_s1, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_clock_crossing_master_ddr2_s1_module burstcount_fifo_for_clock_crossing_master_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (clock_crossing_master_ddr2_s1_selected_burstcount),
      .data_out             (clock_crossing_master_ddr2_s1_transaction_burst_count),
      .empty                (clock_crossing_master_ddr2_s1_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read & clock_crossing_master_ddr2_s1_load_fifo & ~(clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst & clock_crossing_master_ddr2_s1_burstcount_fifo_empty))
    );

  //clock_crossing_master_ddr2_s1 current burst minus one, which is an e_assign
  assign clock_crossing_master_ddr2_s1_current_burst_minus_one = clock_crossing_master_ddr2_s1_current_burst - 1;

  //what to load in current_burst, for clock_crossing_master_ddr2_s1, which is an e_mux
  assign clock_crossing_master_ddr2_s1_next_burst_count = (((in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read) & ~clock_crossing_master_ddr2_s1_load_fifo))? clock_crossing_master_ddr2_s1_selected_burstcount :
    ((in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read & clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst & clock_crossing_master_ddr2_s1_burstcount_fifo_empty))? clock_crossing_master_ddr2_s1_selected_burstcount :
    (clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst)? clock_crossing_master_ddr2_s1_transaction_burst_count :
    clock_crossing_master_ddr2_s1_current_burst_minus_one;

  //the current burst count for clock_crossing_master_ddr2_s1, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_current_burst <= 0;
      else if (clock_crossing_master_ddr2_s1_readdatavalid_from_sa | (~clock_crossing_master_ddr2_s1_load_fifo & (in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read)))
          clock_crossing_master_ddr2_s1_current_burst <= clock_crossing_master_ddr2_s1_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_clock_crossing_master_ddr2_s1_load_fifo = (~clock_crossing_master_ddr2_s1_load_fifo)? 1 :
    (((in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read) & clock_crossing_master_ddr2_s1_load_fifo))? 1 :
    ~clock_crossing_master_ddr2_s1_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_load_fifo <= 0;
      else if ((in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read) & ~clock_crossing_master_ddr2_s1_load_fifo | clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst)
          clock_crossing_master_ddr2_s1_load_fifo <= p0_clock_crossing_master_ddr2_s1_load_fifo;
    end


  //the last cycle in the burst for clock_crossing_master_ddr2_s1, which is an e_assign
  assign clock_crossing_master_ddr2_s1_this_cycle_is_the_last_burst = ~(|clock_crossing_master_ddr2_s1_current_burst_minus_one) & clock_crossing_master_ddr2_s1_readdatavalid_from_sa;

  //rdv_fifo_for_master_read_avalon_master_to_clock_crossing_master_ddr2_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_master_read_avalon_master_to_clock_crossing_master_ddr2_s1_module rdv_fifo_for_master_read_avalon_master_to_clock_crossing_master_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (master_read_granted_clock_crossing_master_ddr2_s1),
      .data_out             (master_read_rdv_fifo_output_from_clock_crossing_master_ddr2_s1),
      .empty                (),
      .fifo_contains_ones_n (master_read_rdv_fifo_empty_clock_crossing_master_ddr2_s1),
      .full                 (),
      .read                 (clock_crossing_master_ddr2_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_master_ddr2_s1_waits_for_read)
    );

  assign master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register = ~master_read_rdv_fifo_empty_clock_crossing_master_ddr2_s1;
  //local readdatavalid master_read_read_data_valid_clock_crossing_master_ddr2_s1, which is an e_mux
  assign master_read_read_data_valid_clock_crossing_master_ddr2_s1 = (clock_crossing_master_ddr2_s1_readdatavalid_from_sa & master_read_rdv_fifo_output_from_clock_crossing_master_ddr2_s1) & ~ master_read_rdv_fifo_empty_clock_crossing_master_ddr2_s1;

  //assign clock_crossing_master_ddr2_s1_endofpacket_from_sa = clock_crossing_master_ddr2_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_master_ddr2_s1_endofpacket_from_sa = clock_crossing_master_ddr2_s1_endofpacket;

  assign master_write_requests_clock_crossing_master_ddr2_s1 = ((1) & (master_write_avalon_master_write)) & master_write_avalon_master_write;
  //master_read/avalon_master granted clock_crossing_master_ddr2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_master_read_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 <= 0;
      else 
        last_cycle_master_read_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 <= master_read_saved_grant_clock_crossing_master_ddr2_s1 ? 1 : (clock_crossing_master_ddr2_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_master_read_avalon_master_granted_slave_clock_crossing_master_ddr2_s1;
    end


  //master_read_avalon_master_continuerequest continued request, which is an e_mux
  assign master_read_avalon_master_continuerequest = last_cycle_master_read_avalon_master_granted_slave_clock_crossing_master_ddr2_s1 & 1;

  assign master_write_qualified_request_clock_crossing_master_ddr2_s1 = master_write_requests_clock_crossing_master_ddr2_s1 & ~(master_read_avalon_master_arbiterlock);
  //clock_crossing_master_ddr2_s1_writedata mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_writedata = master_write_avalon_master_writedata;

  //allow new arb cycle for clock_crossing_master_ddr2/s1, which is an e_assign
  assign clock_crossing_master_ddr2_s1_allow_new_arb_cycle = ~master_read_avalon_master_arbiterlock & ~master_write_avalon_master_arbiterlock;

  //master_write/avalon_master assignment into master qualified-requests vector for clock_crossing_master_ddr2/s1, which is an e_assign
  assign clock_crossing_master_ddr2_s1_master_qreq_vector[0] = master_write_qualified_request_clock_crossing_master_ddr2_s1;

  //master_write/avalon_master grant clock_crossing_master_ddr2/s1, which is an e_assign
  assign master_write_granted_clock_crossing_master_ddr2_s1 = clock_crossing_master_ddr2_s1_grant_vector[0];

  //master_write/avalon_master saved-grant clock_crossing_master_ddr2/s1, which is an e_assign
  assign master_write_saved_grant_clock_crossing_master_ddr2_s1 = clock_crossing_master_ddr2_s1_arb_winner[0];

  //master_read/avalon_master assignment into master qualified-requests vector for clock_crossing_master_ddr2/s1, which is an e_assign
  assign clock_crossing_master_ddr2_s1_master_qreq_vector[1] = master_read_qualified_request_clock_crossing_master_ddr2_s1;

  //master_read/avalon_master grant clock_crossing_master_ddr2/s1, which is an e_assign
  assign master_read_granted_clock_crossing_master_ddr2_s1 = clock_crossing_master_ddr2_s1_grant_vector[1];

  //master_read/avalon_master saved-grant clock_crossing_master_ddr2/s1, which is an e_assign
  assign master_read_saved_grant_clock_crossing_master_ddr2_s1 = clock_crossing_master_ddr2_s1_arb_winner[1];

  //clock_crossing_master_ddr2/s1 chosen-master double-vector, which is an e_assign
  assign clock_crossing_master_ddr2_s1_chosen_master_double_vector = {clock_crossing_master_ddr2_s1_master_qreq_vector, clock_crossing_master_ddr2_s1_master_qreq_vector} & ({~clock_crossing_master_ddr2_s1_master_qreq_vector, ~clock_crossing_master_ddr2_s1_master_qreq_vector} + clock_crossing_master_ddr2_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign clock_crossing_master_ddr2_s1_arb_winner = (clock_crossing_master_ddr2_s1_allow_new_arb_cycle & | clock_crossing_master_ddr2_s1_grant_vector) ? clock_crossing_master_ddr2_s1_grant_vector : clock_crossing_master_ddr2_s1_saved_chosen_master_vector;

  //saved clock_crossing_master_ddr2_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_saved_chosen_master_vector <= 0;
      else if (clock_crossing_master_ddr2_s1_allow_new_arb_cycle)
          clock_crossing_master_ddr2_s1_saved_chosen_master_vector <= |clock_crossing_master_ddr2_s1_grant_vector ? clock_crossing_master_ddr2_s1_grant_vector : clock_crossing_master_ddr2_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign clock_crossing_master_ddr2_s1_grant_vector = {(clock_crossing_master_ddr2_s1_chosen_master_double_vector[1] | clock_crossing_master_ddr2_s1_chosen_master_double_vector[3]),
    (clock_crossing_master_ddr2_s1_chosen_master_double_vector[0] | clock_crossing_master_ddr2_s1_chosen_master_double_vector[2])};

  //clock_crossing_master_ddr2/s1 chosen master rotated left, which is an e_assign
  assign clock_crossing_master_ddr2_s1_chosen_master_rot_left = (clock_crossing_master_ddr2_s1_arb_winner << 1) ? (clock_crossing_master_ddr2_s1_arb_winner << 1) : 1;

  //clock_crossing_master_ddr2/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_arb_addend <= 1;
      else if (|clock_crossing_master_ddr2_s1_grant_vector)
          clock_crossing_master_ddr2_s1_arb_addend <= clock_crossing_master_ddr2_s1_end_xfer? clock_crossing_master_ddr2_s1_chosen_master_rot_left : clock_crossing_master_ddr2_s1_grant_vector;
    end


  //clock_crossing_master_ddr2_s1_reset_n assignment, which is an e_assign
  assign clock_crossing_master_ddr2_s1_reset_n = reset_n;

  //clock_crossing_master_ddr2_s1_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_master_ddr2_s1_firsttransfer = clock_crossing_master_ddr2_s1_begins_xfer ? clock_crossing_master_ddr2_s1_unreg_firsttransfer : clock_crossing_master_ddr2_s1_reg_firsttransfer;

  //clock_crossing_master_ddr2_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_master_ddr2_s1_unreg_firsttransfer = ~(clock_crossing_master_ddr2_s1_slavearbiterlockenable & clock_crossing_master_ddr2_s1_any_continuerequest);

  //clock_crossing_master_ddr2_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_reg_firsttransfer <= 1'b1;
      else if (clock_crossing_master_ddr2_s1_begins_xfer)
          clock_crossing_master_ddr2_s1_reg_firsttransfer <= clock_crossing_master_ddr2_s1_unreg_firsttransfer;
    end


  //clock_crossing_master_ddr2_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign clock_crossing_master_ddr2_s1_next_bbt_burstcount = ((((clock_crossing_master_ddr2_s1_write) && (clock_crossing_master_ddr2_s1_bbt_burstcounter == 0))))? (clock_crossing_master_ddr2_s1_burstcount - 1) :
    ((((clock_crossing_master_ddr2_s1_read) && (clock_crossing_master_ddr2_s1_bbt_burstcounter == 0))))? 0 :
    (clock_crossing_master_ddr2_s1_bbt_burstcounter - 1);

  //clock_crossing_master_ddr2_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_s1_bbt_burstcounter <= 0;
      else if (clock_crossing_master_ddr2_s1_begins_xfer)
          clock_crossing_master_ddr2_s1_bbt_burstcounter <= clock_crossing_master_ddr2_s1_next_bbt_burstcount;
    end


  //clock_crossing_master_ddr2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign clock_crossing_master_ddr2_s1_beginbursttransfer_internal = clock_crossing_master_ddr2_s1_begins_xfer & (clock_crossing_master_ddr2_s1_bbt_burstcounter == 0);

  //clock_crossing_master_ddr2_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign clock_crossing_master_ddr2_s1_arbitration_holdoff_internal = clock_crossing_master_ddr2_s1_begins_xfer & clock_crossing_master_ddr2_s1_firsttransfer;

  //clock_crossing_master_ddr2_s1_read assignment, which is an e_mux
  assign clock_crossing_master_ddr2_s1_read = master_read_granted_clock_crossing_master_ddr2_s1 & master_read_avalon_master_read;

  //clock_crossing_master_ddr2_s1_write assignment, which is an e_mux
  assign clock_crossing_master_ddr2_s1_write = master_write_granted_clock_crossing_master_ddr2_s1 & master_write_avalon_master_write;

  assign shifted_address_to_clock_crossing_master_ddr2_s1_from_master_read_avalon_master = master_read_avalon_master_address_to_slave;
  //clock_crossing_master_ddr2_s1_address mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_address = (master_read_granted_clock_crossing_master_ddr2_s1)? (shifted_address_to_clock_crossing_master_ddr2_s1_from_master_read_avalon_master >> 5) :
    (shifted_address_to_clock_crossing_master_ddr2_s1_from_master_write_avalon_master >> 5);

  assign shifted_address_to_clock_crossing_master_ddr2_s1_from_master_write_avalon_master = master_write_avalon_master_address_to_slave;
  //slaveid clock_crossing_master_ddr2_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_nativeaddress = (master_read_granted_clock_crossing_master_ddr2_s1)? (master_read_avalon_master_address_to_slave >> 5) :
    (master_write_avalon_master_address_to_slave >> 5);

  //d1_clock_crossing_master_ddr2_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_clock_crossing_master_ddr2_s1_end_xfer <= 1;
      else 
        d1_clock_crossing_master_ddr2_s1_end_xfer <= clock_crossing_master_ddr2_s1_end_xfer;
    end


  //clock_crossing_master_ddr2_s1_waits_for_read in a cycle, which is an e_mux
  assign clock_crossing_master_ddr2_s1_waits_for_read = clock_crossing_master_ddr2_s1_in_a_read_cycle & clock_crossing_master_ddr2_s1_waitrequest_from_sa;

  //clock_crossing_master_ddr2_s1_in_a_read_cycle assignment, which is an e_assign
  assign clock_crossing_master_ddr2_s1_in_a_read_cycle = master_read_granted_clock_crossing_master_ddr2_s1 & master_read_avalon_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = clock_crossing_master_ddr2_s1_in_a_read_cycle;

  //clock_crossing_master_ddr2_s1_waits_for_write in a cycle, which is an e_mux
  assign clock_crossing_master_ddr2_s1_waits_for_write = clock_crossing_master_ddr2_s1_in_a_write_cycle & clock_crossing_master_ddr2_s1_waitrequest_from_sa;

  //clock_crossing_master_ddr2_s1_in_a_write_cycle assignment, which is an e_assign
  assign clock_crossing_master_ddr2_s1_in_a_write_cycle = master_write_granted_clock_crossing_master_ddr2_s1 & master_write_avalon_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = clock_crossing_master_ddr2_s1_in_a_write_cycle;

  assign wait_for_clock_crossing_master_ddr2_s1_counter = 0;
  //clock_crossing_master_ddr2_s1_byteenable byte enable port mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_byteenable = (master_write_granted_clock_crossing_master_ddr2_s1)? master_write_avalon_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign clock_crossing_master_ddr2_s1_burstcount = (master_read_granted_clock_crossing_master_ddr2_s1)? master_read_avalon_master_burstcount :
    (master_write_granted_clock_crossing_master_ddr2_s1)? master_write_avalon_master_burstcount :
    1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_master_ddr2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //master_read/avalon_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (master_read_requests_clock_crossing_master_ddr2_s1 && (master_read_avalon_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: master_read/avalon_master drove 0 on its 'burstcount' port while accessing slave clock_crossing_master_ddr2/s1", $time);
          $stop;
        end
    end


  //master_write/avalon_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (master_write_requests_clock_crossing_master_ddr2_s1 && (master_write_avalon_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: master_write/avalon_master drove 0 on its 'burstcount' port while accessing slave clock_crossing_master_ddr2/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (master_read_granted_clock_crossing_master_ddr2_s1 + master_write_granted_clock_crossing_master_ddr2_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (master_read_saved_grant_clock_crossing_master_ddr2_s1 + master_write_saved_grant_clock_crossing_master_ddr2_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_master_ddr2_m1_arbitrator (
                                                  // inputs:
                                                   SS_OCT_SOPC_burst_0_upstream_readdata_from_sa,
                                                   SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa,
                                                   clk,
                                                   clock_crossing_master_ddr2_m1_address,
                                                   clock_crossing_master_ddr2_m1_burstcount,
                                                   clock_crossing_master_ddr2_m1_byteenable,
                                                   clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream,
                                                   clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream,
                                                   clock_crossing_master_ddr2_m1_read,
                                                   clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream,
                                                   clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register,
                                                   clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream,
                                                   clock_crossing_master_ddr2_m1_write,
                                                   clock_crossing_master_ddr2_m1_writedata,
                                                   d1_SS_OCT_SOPC_burst_0_upstream_end_xfer,
                                                   reset_n,

                                                  // outputs:
                                                   clock_crossing_master_ddr2_m1_address_to_slave,
                                                   clock_crossing_master_ddr2_m1_latency_counter,
                                                   clock_crossing_master_ddr2_m1_readdata,
                                                   clock_crossing_master_ddr2_m1_readdatavalid,
                                                   clock_crossing_master_ddr2_m1_reset_n,
                                                   clock_crossing_master_ddr2_m1_waitrequest
                                                )
;

  output  [ 29: 0] clock_crossing_master_ddr2_m1_address_to_slave;
  output           clock_crossing_master_ddr2_m1_latency_counter;
  output  [255: 0] clock_crossing_master_ddr2_m1_readdata;
  output           clock_crossing_master_ddr2_m1_readdatavalid;
  output           clock_crossing_master_ddr2_m1_reset_n;
  output           clock_crossing_master_ddr2_m1_waitrequest;
  input   [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata_from_sa;
  input            SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;
  input            clk;
  input   [ 29: 0] clock_crossing_master_ddr2_m1_address;
  input   [  3: 0] clock_crossing_master_ddr2_m1_burstcount;
  input   [ 31: 0] clock_crossing_master_ddr2_m1_byteenable;
  input            clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream;
  input            clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream;
  input            clock_crossing_master_ddr2_m1_read;
  input            clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream;
  input            clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register;
  input            clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream;
  input            clock_crossing_master_ddr2_m1_write;
  input   [255: 0] clock_crossing_master_ddr2_m1_writedata;
  input            d1_SS_OCT_SOPC_burst_0_upstream_end_xfer;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 29: 0] clock_crossing_master_ddr2_m1_address_last_time;
  wire    [ 29: 0] clock_crossing_master_ddr2_m1_address_to_slave;
  reg     [  3: 0] clock_crossing_master_ddr2_m1_burstcount_last_time;
  reg     [ 31: 0] clock_crossing_master_ddr2_m1_byteenable_last_time;
  wire             clock_crossing_master_ddr2_m1_latency_counter;
  reg              clock_crossing_master_ddr2_m1_read_last_time;
  wire    [255: 0] clock_crossing_master_ddr2_m1_readdata;
  wire             clock_crossing_master_ddr2_m1_readdatavalid;
  wire             clock_crossing_master_ddr2_m1_reset_n;
  wire             clock_crossing_master_ddr2_m1_run;
  wire             clock_crossing_master_ddr2_m1_waitrequest;
  reg              clock_crossing_master_ddr2_m1_write_last_time;
  reg     [255: 0] clock_crossing_master_ddr2_m1_writedata_last_time;
  wire             pre_flush_clock_crossing_master_ddr2_m1_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream | ~clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream) & ((~clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream | ~(clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write) | (1 & ~SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa & (clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write)))) & ((~clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream | ~(clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write) | (1 & ~SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa & (clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write))));

  //cascaded wait assignment, which is an e_assign
  assign clock_crossing_master_ddr2_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign clock_crossing_master_ddr2_m1_address_to_slave = clock_crossing_master_ddr2_m1_address[29 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_clock_crossing_master_ddr2_m1_readdatavalid = clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign clock_crossing_master_ddr2_m1_readdatavalid = 0 |
    pre_flush_clock_crossing_master_ddr2_m1_readdatavalid;

  //clock_crossing_master_ddr2/m1 readdata mux, which is an e_mux
  assign clock_crossing_master_ddr2_m1_readdata = SS_OCT_SOPC_burst_0_upstream_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign clock_crossing_master_ddr2_m1_waitrequest = ~clock_crossing_master_ddr2_m1_run;

  //latent max counter, which is an e_assign
  assign clock_crossing_master_ddr2_m1_latency_counter = 0;

  //clock_crossing_master_ddr2_m1_reset_n assignment, which is an e_assign
  assign clock_crossing_master_ddr2_m1_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_master_ddr2_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_address_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_address_last_time <= clock_crossing_master_ddr2_m1_address;
    end


  //clock_crossing_master_ddr2/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= clock_crossing_master_ddr2_m1_waitrequest & (clock_crossing_master_ddr2_m1_read | clock_crossing_master_ddr2_m1_write);
    end


  //clock_crossing_master_ddr2_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_address != clock_crossing_master_ddr2_m1_address_last_time))
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_master_ddr2_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_burstcount_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_burstcount_last_time <= clock_crossing_master_ddr2_m1_burstcount;
    end


  //clock_crossing_master_ddr2_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_burstcount != clock_crossing_master_ddr2_m1_burstcount_last_time))
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_master_ddr2_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_byteenable_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_byteenable_last_time <= clock_crossing_master_ddr2_m1_byteenable;
    end


  //clock_crossing_master_ddr2_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_byteenable != clock_crossing_master_ddr2_m1_byteenable_last_time))
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_master_ddr2_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_read_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_read_last_time <= clock_crossing_master_ddr2_m1_read;
    end


  //clock_crossing_master_ddr2_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_read != clock_crossing_master_ddr2_m1_read_last_time))
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_master_ddr2_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_write_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_write_last_time <= clock_crossing_master_ddr2_m1_write;
    end


  //clock_crossing_master_ddr2_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_write != clock_crossing_master_ddr2_m1_write_last_time))
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_master_ddr2_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_master_ddr2_m1_writedata_last_time <= 0;
      else 
        clock_crossing_master_ddr2_m1_writedata_last_time <= clock_crossing_master_ddr2_m1_writedata;
    end


  //clock_crossing_master_ddr2_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_master_ddr2_m1_writedata != clock_crossing_master_ddr2_m1_writedata_last_time) & clock_crossing_master_ddr2_m1_write)
        begin
          $write("%0d ns: clock_crossing_master_ddr2_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_master_ddr2_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_data_master_address_to_slave,
                                           cpu_data_master_byteenable,
                                           cpu_data_master_debugaccess,
                                           cpu_data_master_latency_counter,
                                           cpu_data_master_read,
                                           cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                           cpu_data_master_write,
                                           cpu_data_master_writedata,
                                           cpu_instruction_master_address_to_slave,
                                           cpu_instruction_master_latency_counter,
                                           cpu_instruction_master_read,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           reset_n,

                                          // outputs:
                                           cpu_data_master_granted_cpu_jtag_debug_module,
                                           cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_data_master_requests_cpu_jtag_debug_module,
                                           cpu_instruction_master_granted_cpu_jtag_debug_module,
                                           cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_instruction_master_requests_cpu_jtag_debug_module,
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer
                                        )
;

  output           cpu_data_master_granted_cpu_jtag_debug_module;
  output           cpu_data_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_data_master_requests_cpu_jtag_debug_module;
  output           cpu_instruction_master_granted_cpu_jtag_debug_module;
  output           cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_instruction_master_requests_cpu_jtag_debug_module;
  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 30: 0] cpu_instruction_master_address_to_slave;
  input   [  1: 0] cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_saved_grant_cpu_jtag_debug_module;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_saved_grant_cpu_jtag_debug_module;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_jtag_debug_module_arb_addend;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg     [  1: 0] cpu_jtag_debug_module_arb_share_counter;
  wire    [  1: 0] cpu_jtag_debug_module_arb_share_counter_next_value;
  wire    [  1: 0] cpu_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_jtag_debug_module_arb_winner;
  wire             cpu_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
  reg              last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
  wire    [ 30: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master;
  wire    [ 30: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_cpu_jtag_debug_module | cpu_instruction_master_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign cpu_data_master_requests_cpu_jtag_debug_module = ({cpu_data_master_address_to_slave[30 : 11] , 11'b0} == 31'h48111000) & (cpu_data_master_read | cpu_data_master_write);
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module |
    cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector);

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu/data_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_data_master_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //cpu/data_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= cpu_instruction_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_instruction_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module & cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_jtag_debug_module_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_cpu_jtag_debug_module = cpu_data_master_requests_cpu_jtag_debug_module & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //local readdatavalid cpu_data_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_data_master_read_data_valid_cpu_jtag_debug_module = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = cpu_data_master_writedata;

  assign cpu_instruction_master_requests_cpu_jtag_debug_module = (({cpu_instruction_master_address_to_slave[30 : 11] , 11'b0} == 31'h48111000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= cpu_data_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_data_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module & cpu_data_master_requests_cpu_jtag_debug_module;

  assign cpu_instruction_master_qualified_request_cpu_jtag_debug_module = cpu_instruction_master_requests_cpu_jtag_debug_module & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0))) | cpu_data_master_arbiterlock);
  //local readdatavalid cpu_instruction_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_instruction_master_read_data_valid_cpu_jtag_debug_module = cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[0] = cpu_instruction_master_qualified_request_cpu_jtag_debug_module;

  //cpu/instruction_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[0];

  //cpu/instruction_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[0] && cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu/data_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[1] = cpu_data_master_qualified_request_cpu_jtag_debug_module;

  //cpu/data_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[1];

  //cpu/data_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[1] && cpu_data_master_requests_cpu_jtag_debug_module;

  //cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_double_vector = {cpu_jtag_debug_module_master_qreq_vector, cpu_jtag_debug_module_master_qreq_vector} & ({~cpu_jtag_debug_module_master_qreq_vector, ~cpu_jtag_debug_module_master_qreq_vector} + cpu_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_jtag_debug_module_arb_winner = (cpu_jtag_debug_module_allow_new_arb_cycle & | cpu_jtag_debug_module_grant_vector) ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_jtag_debug_module_allow_new_arb_cycle)
          cpu_jtag_debug_module_saved_chosen_master_vector <= |cpu_jtag_debug_module_grant_vector ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_jtag_debug_module_grant_vector = {(cpu_jtag_debug_module_chosen_master_double_vector[1] | cpu_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_jtag_debug_module_chosen_master_double_vector[0] | cpu_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_rot_left = (cpu_jtag_debug_module_arb_winner << 1) ? (cpu_jtag_debug_module_arb_winner << 1) : 1;

  //cpu/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_jtag_debug_module_grant_vector)
          cpu_jtag_debug_module_arb_addend <= cpu_jtag_debug_module_end_xfer? cpu_jtag_debug_module_chosen_master_rot_left : cpu_jtag_debug_module_grant_vector;
    end


  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = cpu_data_master_granted_cpu_jtag_debug_module | cpu_instruction_master_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_jtag_debug_module_arbitration_holdoff_internal = cpu_jtag_debug_module_begins_xfer & cpu_jtag_debug_module_firsttransfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master = cpu_data_master_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = (cpu_data_master_granted_cpu_jtag_debug_module)? (shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master >> 2) :
    (shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master >> 2);

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = (cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_cpu_jtag_debug_module + cpu_instruction_master_granted_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_cpu_jtag_debug_module + cpu_instruction_master_saved_grant_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     SS_OCT_SOPC_clock_0_in_readdata_from_sa,
                                     SS_OCT_SOPC_clock_0_in_waitrequest_from_sa,
                                     clk,
                                     clock_crossing_ddr2_cpu_s1_readdata_from_sa,
                                     clock_crossing_ddr2_cpu_s1_waitrequest_from_sa,
                                     cpu_data_master_address,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_byteenable_ext_flash_s1,
                                     cpu_data_master_granted_SS_OCT_SOPC_clock_0_in,
                                     cpu_data_master_granted_clock_crossing_ddr2_cpu_s1,
                                     cpu_data_master_granted_cpu_jtag_debug_module,
                                     cpu_data_master_granted_descriptor_memory_s1,
                                     cpu_data_master_granted_ext_flash_s1,
                                     cpu_data_master_granted_high_res_timer_s1,
                                     cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_granted_onchip_memory_s1,
                                     cpu_data_master_granted_packet_memory_s1,
                                     cpu_data_master_granted_sgdma_rx_csr,
                                     cpu_data_master_granted_sgdma_tx_csr,
                                     cpu_data_master_granted_sys_timer_s1,
                                     cpu_data_master_granted_sysid_control_slave,
                                     cpu_data_master_granted_tse_mac_control_port,
                                     cpu_data_master_granted_vol_recording_done_pio_s1,
                                     cpu_data_master_granted_vol_transfer_done_pio_s1,
                                     cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in,
                                     cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1,
                                     cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                     cpu_data_master_qualified_request_descriptor_memory_s1,
                                     cpu_data_master_qualified_request_ext_flash_s1,
                                     cpu_data_master_qualified_request_high_res_timer_s1,
                                     cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_qualified_request_onchip_memory_s1,
                                     cpu_data_master_qualified_request_packet_memory_s1,
                                     cpu_data_master_qualified_request_sgdma_rx_csr,
                                     cpu_data_master_qualified_request_sgdma_tx_csr,
                                     cpu_data_master_qualified_request_sys_timer_s1,
                                     cpu_data_master_qualified_request_sysid_control_slave,
                                     cpu_data_master_qualified_request_tse_mac_control_port,
                                     cpu_data_master_qualified_request_vol_recording_done_pio_s1,
                                     cpu_data_master_qualified_request_vol_transfer_done_pio_s1,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in,
                                     cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1,
                                     cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                     cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                     cpu_data_master_read_data_valid_descriptor_memory_s1,
                                     cpu_data_master_read_data_valid_ext_flash_s1,
                                     cpu_data_master_read_data_valid_high_res_timer_s1,
                                     cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_read_data_valid_onchip_memory_s1,
                                     cpu_data_master_read_data_valid_packet_memory_s1,
                                     cpu_data_master_read_data_valid_sgdma_rx_csr,
                                     cpu_data_master_read_data_valid_sgdma_tx_csr,
                                     cpu_data_master_read_data_valid_sys_timer_s1,
                                     cpu_data_master_read_data_valid_sysid_control_slave,
                                     cpu_data_master_read_data_valid_tse_mac_control_port,
                                     cpu_data_master_read_data_valid_vol_recording_done_pio_s1,
                                     cpu_data_master_read_data_valid_vol_transfer_done_pio_s1,
                                     cpu_data_master_requests_SS_OCT_SOPC_clock_0_in,
                                     cpu_data_master_requests_clock_crossing_ddr2_cpu_s1,
                                     cpu_data_master_requests_cpu_jtag_debug_module,
                                     cpu_data_master_requests_descriptor_memory_s1,
                                     cpu_data_master_requests_ext_flash_s1,
                                     cpu_data_master_requests_high_res_timer_s1,
                                     cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
                                     cpu_data_master_requests_onchip_memory_s1,
                                     cpu_data_master_requests_packet_memory_s1,
                                     cpu_data_master_requests_sgdma_rx_csr,
                                     cpu_data_master_requests_sgdma_tx_csr,
                                     cpu_data_master_requests_sys_timer_s1,
                                     cpu_data_master_requests_sysid_control_slave,
                                     cpu_data_master_requests_tse_mac_control_port,
                                     cpu_data_master_requests_vol_recording_done_pio_s1,
                                     cpu_data_master_requests_vol_transfer_done_pio_s1,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     cpu_jtag_debug_module_readdata_from_sa,
                                     d1_SS_OCT_SOPC_clock_0_in_end_xfer,
                                     d1_clock_crossing_ddr2_cpu_s1_end_xfer,
                                     d1_cpu_jtag_debug_module_end_xfer,
                                     d1_descriptor_memory_s1_end_xfer,
                                     d1_flash_tristate_bridge_avalon_slave_end_xfer,
                                     d1_high_res_timer_s1_end_xfer,
                                     d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                     d1_onchip_memory_s1_end_xfer,
                                     d1_packet_memory_s1_end_xfer,
                                     d1_sgdma_rx_csr_end_xfer,
                                     d1_sgdma_tx_csr_end_xfer,
                                     d1_sys_timer_s1_end_xfer,
                                     d1_sysid_control_slave_end_xfer,
                                     d1_tse_mac_control_port_end_xfer,
                                     d1_vol_recording_done_pio_s1_end_xfer,
                                     d1_vol_transfer_done_pio_s1_end_xfer,
                                     descriptor_memory_s1_readdata_from_sa,
                                     ext_flash_s1_wait_counter_eq_0,
                                     high_res_timer_s1_irq_from_sa,
                                     high_res_timer_s1_readdata_from_sa,
                                     incoming_flash_tristate_bridge_data_with_Xs_converted_to_0,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                     jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                     onchip_memory_s1_readdata_from_sa,
                                     packet_memory_s1_readdata_from_sa,
                                     reset_n,
                                     sgdma_rx_csr_irq_from_sa,
                                     sgdma_rx_csr_readdata_from_sa,
                                     sgdma_tx_csr_irq_from_sa,
                                     sgdma_tx_csr_readdata_from_sa,
                                     sys_timer_s1_irq_from_sa,
                                     sys_timer_s1_readdata_from_sa,
                                     sysid_control_slave_readdata_from_sa,
                                     tse_mac_control_port_readdata_from_sa,
                                     tse_mac_control_port_waitrequest_from_sa,
                                     vol_recording_done_pio_s1_readdata_from_sa,
                                     vol_transfer_done_pio_s1_readdata_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_dbs_address,
                                     cpu_data_master_dbs_write_16,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 30: 0] cpu_data_master_address_to_slave;
  output  [  1: 0] cpu_data_master_dbs_address;
  output  [ 15: 0] cpu_data_master_dbs_write_16;
  output  [ 31: 0] cpu_data_master_irq;
  output  [  1: 0] cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input   [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata_from_sa;
  input            SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;
  input            clk;
  input   [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata_from_sa;
  input            clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;
  input   [ 30: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_byteenable_ext_flash_s1;
  input            cpu_data_master_granted_SS_OCT_SOPC_clock_0_in;
  input            cpu_data_master_granted_clock_crossing_ddr2_cpu_s1;
  input            cpu_data_master_granted_cpu_jtag_debug_module;
  input            cpu_data_master_granted_descriptor_memory_s1;
  input            cpu_data_master_granted_ext_flash_s1;
  input            cpu_data_master_granted_high_res_timer_s1;
  input            cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_granted_onchip_memory_s1;
  input            cpu_data_master_granted_packet_memory_s1;
  input            cpu_data_master_granted_sgdma_rx_csr;
  input            cpu_data_master_granted_sgdma_tx_csr;
  input            cpu_data_master_granted_sys_timer_s1;
  input            cpu_data_master_granted_sysid_control_slave;
  input            cpu_data_master_granted_tse_mac_control_port;
  input            cpu_data_master_granted_vol_recording_done_pio_s1;
  input            cpu_data_master_granted_vol_transfer_done_pio_s1;
  input            cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in;
  input            cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1;
  input            cpu_data_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_data_master_qualified_request_descriptor_memory_s1;
  input            cpu_data_master_qualified_request_ext_flash_s1;
  input            cpu_data_master_qualified_request_high_res_timer_s1;
  input            cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_qualified_request_onchip_memory_s1;
  input            cpu_data_master_qualified_request_packet_memory_s1;
  input            cpu_data_master_qualified_request_sgdma_rx_csr;
  input            cpu_data_master_qualified_request_sgdma_tx_csr;
  input            cpu_data_master_qualified_request_sys_timer_s1;
  input            cpu_data_master_qualified_request_sysid_control_slave;
  input            cpu_data_master_qualified_request_tse_mac_control_port;
  input            cpu_data_master_qualified_request_vol_recording_done_pio_s1;
  input            cpu_data_master_qualified_request_vol_transfer_done_pio_s1;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_data_master_read_data_valid_descriptor_memory_s1;
  input            cpu_data_master_read_data_valid_ext_flash_s1;
  input            cpu_data_master_read_data_valid_high_res_timer_s1;
  input            cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_read_data_valid_onchip_memory_s1;
  input            cpu_data_master_read_data_valid_packet_memory_s1;
  input            cpu_data_master_read_data_valid_sgdma_rx_csr;
  input            cpu_data_master_read_data_valid_sgdma_tx_csr;
  input            cpu_data_master_read_data_valid_sys_timer_s1;
  input            cpu_data_master_read_data_valid_sysid_control_slave;
  input            cpu_data_master_read_data_valid_tse_mac_control_port;
  input            cpu_data_master_read_data_valid_vol_recording_done_pio_s1;
  input            cpu_data_master_read_data_valid_vol_transfer_done_pio_s1;
  input            cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;
  input            cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;
  input            cpu_data_master_requests_cpu_jtag_debug_module;
  input            cpu_data_master_requests_descriptor_memory_s1;
  input            cpu_data_master_requests_ext_flash_s1;
  input            cpu_data_master_requests_high_res_timer_s1;
  input            cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  input            cpu_data_master_requests_onchip_memory_s1;
  input            cpu_data_master_requests_packet_memory_s1;
  input            cpu_data_master_requests_sgdma_rx_csr;
  input            cpu_data_master_requests_sgdma_tx_csr;
  input            cpu_data_master_requests_sys_timer_s1;
  input            cpu_data_master_requests_sysid_control_slave;
  input            cpu_data_master_requests_tse_mac_control_port;
  input            cpu_data_master_requests_vol_recording_done_pio_s1;
  input            cpu_data_master_requests_vol_transfer_done_pio_s1;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_SS_OCT_SOPC_clock_0_in_end_xfer;
  input            d1_clock_crossing_ddr2_cpu_s1_end_xfer;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_descriptor_memory_s1_end_xfer;
  input            d1_flash_tristate_bridge_avalon_slave_end_xfer;
  input            d1_high_res_timer_s1_end_xfer;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_onchip_memory_s1_end_xfer;
  input            d1_packet_memory_s1_end_xfer;
  input            d1_sgdma_rx_csr_end_xfer;
  input            d1_sgdma_tx_csr_end_xfer;
  input            d1_sys_timer_s1_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_tse_mac_control_port_end_xfer;
  input            d1_vol_recording_done_pio_s1_end_xfer;
  input            d1_vol_transfer_done_pio_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            ext_flash_s1_wait_counter_eq_0;
  input            high_res_timer_s1_irq_from_sa;
  input   [ 15: 0] high_res_timer_s1_readdata_from_sa;
  input   [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory_s1_readdata_from_sa;
  input   [ 31: 0] packet_memory_s1_readdata_from_sa;
  input            reset_n;
  input            sgdma_rx_csr_irq_from_sa;
  input   [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  input            sgdma_tx_csr_irq_from_sa;
  input   [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  input            sys_timer_s1_irq_from_sa;
  input   [ 15: 0] sys_timer_s1_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 31: 0] tse_mac_control_port_readdata_from_sa;
  input            tse_mac_control_port_waitrequest_from_sa;
  input            vol_recording_done_pio_s1_readdata_from_sa;
  input            vol_transfer_done_pio_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 30: 0] cpu_data_master_address_last_time;
  wire    [ 30: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_data_master_dbs_address;
  wire    [  1: 0] cpu_data_master_dbs_increment;
  reg     [  1: 0] cpu_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_data_master_dbs_write_16;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg     [  1: 0] cpu_data_master_latency_counter;
  wire    [  1: 0] cpu_data_master_next_dbs_rdv_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [  1: 0] p1_cpu_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in | ~cpu_data_master_requests_SS_OCT_SOPC_clock_0_in) & ((~cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~SS_OCT_SOPC_clock_0_in_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~SS_OCT_SOPC_clock_0_in_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1 | ~cpu_data_master_requests_clock_crossing_ddr2_cpu_s1) & ((~cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~clock_crossing_ddr2_cpu_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~clock_crossing_ddr2_cpu_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_requests_cpu_jtag_debug_module) & (cpu_data_master_granted_cpu_jtag_debug_module | ~cpu_data_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_descriptor_memory_s1 | ~cpu_data_master_requests_descriptor_memory_s1) & (cpu_data_master_granted_descriptor_memory_s1 | ~cpu_data_master_qualified_request_descriptor_memory_s1) & ((~cpu_data_master_qualified_request_descriptor_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_descriptor_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_ext_flash_s1 | (cpu_data_master_write & !cpu_data_master_byteenable_ext_flash_s1 & cpu_data_master_dbs_address[1]) | ~cpu_data_master_requests_ext_flash_s1);

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_1 & r_2 & r_3;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = (cpu_data_master_granted_ext_flash_s1 | ~cpu_data_master_qualified_request_ext_flash_s1) & ((~cpu_data_master_qualified_request_ext_flash_s1 | ~cpu_data_master_read | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & (cpu_data_master_dbs_address[1]) & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_ext_flash_s1 | ~cpu_data_master_write | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & (cpu_data_master_dbs_address[1]) & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_high_res_timer_s1 | ~cpu_data_master_requests_high_res_timer_s1) & ((~cpu_data_master_qualified_request_high_res_timer_s1 | ~cpu_data_master_read | (1 & ~d1_high_res_timer_s1_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_high_res_timer_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~cpu_data_master_requests_jtag_uart_avalon_jtag_slave) & ((~cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_onchip_memory_s1 | ~cpu_data_master_requests_onchip_memory_s1) & (cpu_data_master_granted_onchip_memory_s1 | ~cpu_data_master_qualified_request_onchip_memory_s1) & ((~cpu_data_master_qualified_request_onchip_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_onchip_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_packet_memory_s1 | ~cpu_data_master_requests_packet_memory_s1) & ((~cpu_data_master_qualified_request_packet_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_packet_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write))));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_requests_sgdma_rx_csr) & ((~cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_read | (1 & ~d1_sgdma_rx_csr_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_requests_sgdma_tx_csr) & ((~cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_read | (1 & ~d1_sgdma_tx_csr_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_sys_timer_s1 | ~cpu_data_master_requests_sys_timer_s1) & ((~cpu_data_master_qualified_request_sys_timer_s1 | ~cpu_data_master_read | (1 & ~d1_sys_timer_s1_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sys_timer_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_sysid_control_slave | ~cpu_data_master_requests_sysid_control_slave) & ((~cpu_data_master_qualified_request_sysid_control_slave | ~cpu_data_master_read | (1 & ~d1_sysid_control_slave_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sysid_control_slave | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_tse_mac_control_port | ~cpu_data_master_requests_tse_mac_control_port) & ((~cpu_data_master_qualified_request_tse_mac_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~tse_mac_control_port_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_tse_mac_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~tse_mac_control_port_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_data_master_qualified_request_vol_recording_done_pio_s1 | ~cpu_data_master_requests_vol_recording_done_pio_s1) & ((~cpu_data_master_qualified_request_vol_recording_done_pio_s1 | ~cpu_data_master_read | (1 & ~d1_vol_recording_done_pio_s1_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_vol_recording_done_pio_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_vol_transfer_done_pio_s1 | ~cpu_data_master_requests_vol_transfer_done_pio_s1) & ((~cpu_data_master_qualified_request_vol_transfer_done_pio_s1 | ~cpu_data_master_read | (1 & ~d1_vol_transfer_done_pio_s1_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_vol_transfer_done_pio_s1 | ~cpu_data_master_write | (1 & cpu_data_master_write)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[30 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_SS_OCT_SOPC_clock_0_in |
    cpu_data_master_granted_clock_crossing_ddr2_cpu_s1 |
    cpu_data_master_granted_cpu_jtag_debug_module |
    cpu_data_master_granted_descriptor_memory_s1 |
    cpu_data_master_granted_ext_flash_s1 |
    cpu_data_master_granted_high_res_timer_s1 |
    cpu_data_master_granted_jtag_uart_avalon_jtag_slave |
    cpu_data_master_granted_onchip_memory_s1 |
    cpu_data_master_granted_packet_memory_s1 |
    cpu_data_master_granted_sgdma_rx_csr |
    cpu_data_master_granted_sgdma_tx_csr |
    cpu_data_master_granted_sys_timer_s1 |
    cpu_data_master_granted_sysid_control_slave |
    cpu_data_master_granted_tse_mac_control_port |
    cpu_data_master_granted_vol_recording_done_pio_s1 |
    cpu_data_master_granted_vol_transfer_done_pio_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1 |
    cpu_data_master_read_data_valid_descriptor_memory_s1 |
    (cpu_data_master_read_data_valid_ext_flash_s1 & dbs_rdv_counter_overflow) |
    cpu_data_master_read_data_valid_onchip_memory_s1 |
    cpu_data_master_read_data_valid_packet_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_cpu_jtag_debug_module |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_high_res_timer_s1 |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sgdma_rx_csr |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sgdma_tx_csr |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sys_timer_s1 |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sysid_control_slave |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_tse_mac_control_port |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_vol_recording_done_pio_s1 |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_vol_transfer_done_pio_s1;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~(cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in & cpu_data_master_read)}} | SS_OCT_SOPC_clock_0_in_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1}} | clock_crossing_ddr2_cpu_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_cpu_jtag_debug_module & cpu_data_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_descriptor_memory_s1}} | descriptor_memory_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_ext_flash_s1}} | {incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_data_master_qualified_request_high_res_timer_s1 & cpu_data_master_read)}} | high_res_timer_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave & cpu_data_master_read)}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_onchip_memory_s1}} | onchip_memory_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_packet_memory_s1}} | packet_memory_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sgdma_rx_csr & cpu_data_master_read)}} | sgdma_rx_csr_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sgdma_tx_csr & cpu_data_master_read)}} | sgdma_tx_csr_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sys_timer_s1 & cpu_data_master_read)}} | sys_timer_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sysid_control_slave & cpu_data_master_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_tse_mac_control_port & cpu_data_master_read)}} | tse_mac_control_port_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_vol_recording_done_pio_s1 & cpu_data_master_read)}} | vol_recording_done_pio_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_vol_transfer_done_pio_s1 & cpu_data_master_read)}} | vol_transfer_done_pio_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else 
        cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {cpu_data_master_requests_descriptor_memory_s1}} & 1) |
    ({2 {cpu_data_master_requests_ext_flash_s1}} & 2) |
    ({2 {cpu_data_master_requests_onchip_memory_s1}} & 1) |
    ({2 {cpu_data_master_requests_packet_memory_s1}} & 1);

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_data_master_requests_ext_flash_s1 & cpu_data_master_write & !cpu_data_master_byteenable_ext_flash_s1)) |
    ((cpu_data_master_granted_ext_flash_s1 & cpu_data_master_read & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer}))) |
    ((cpu_data_master_granted_ext_flash_s1 & cpu_data_master_write & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer})));

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_data_master_dbs_write_16 = (cpu_data_master_dbs_address[1])? cpu_data_master_writedata[31 : 16] :
    cpu_data_master_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign cpu_data_master_dbs_increment = (cpu_data_master_requests_ext_flash_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_data_master_dbs_address + cpu_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_data_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_data_master_next_dbs_rdv_counter = cpu_data_master_dbs_rdv_counter + cpu_data_master_dbs_rdv_counter_inc;

  //cpu_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_data_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_data_master_read_data_valid_ext_flash_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_data_master_dbs_rdv_counter <= cpu_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_data_master_dbs_rdv_counter[1] & ~cpu_data_master_next_dbs_rdv_counter[1];

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    sys_timer_s1_irq_from_sa,
    high_res_timer_s1_irq_from_sa,
    jtag_uart_avalon_jtag_slave_irq_from_sa,
    sgdma_rx_csr_irq_from_sa,
    sgdma_tx_csr_irq_from_sa};


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else 
        cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else 
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else 
        cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else 
        cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else 
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_granted_cpu_jtag_debug_module,
                                            cpu_instruction_master_granted_descriptor_memory_s1,
                                            cpu_instruction_master_granted_ext_flash_s1,
                                            cpu_instruction_master_granted_onchip_memory_s1,
                                            cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                            cpu_instruction_master_qualified_request_descriptor_memory_s1,
                                            cpu_instruction_master_qualified_request_ext_flash_s1,
                                            cpu_instruction_master_qualified_request_onchip_memory_s1,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                            cpu_instruction_master_read_data_valid_descriptor_memory_s1,
                                            cpu_instruction_master_read_data_valid_ext_flash_s1,
                                            cpu_instruction_master_read_data_valid_onchip_memory_s1,
                                            cpu_instruction_master_requests_cpu_jtag_debug_module,
                                            cpu_instruction_master_requests_descriptor_memory_s1,
                                            cpu_instruction_master_requests_ext_flash_s1,
                                            cpu_instruction_master_requests_onchip_memory_s1,
                                            cpu_jtag_debug_module_readdata_from_sa,
                                            d1_cpu_jtag_debug_module_end_xfer,
                                            d1_descriptor_memory_s1_end_xfer,
                                            d1_flash_tristate_bridge_avalon_slave_end_xfer,
                                            d1_onchip_memory_s1_end_xfer,
                                            descriptor_memory_s1_readdata_from_sa,
                                            ext_flash_s1_wait_counter_eq_0,
                                            incoming_flash_tristate_bridge_data,
                                            onchip_memory_s1_readdata_from_sa,
                                            reset_n,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_dbs_address,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 30: 0] cpu_instruction_master_address_to_slave;
  output  [  1: 0] cpu_instruction_master_dbs_address;
  output  [  1: 0] cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 30: 0] cpu_instruction_master_address;
  input            cpu_instruction_master_granted_cpu_jtag_debug_module;
  input            cpu_instruction_master_granted_descriptor_memory_s1;
  input            cpu_instruction_master_granted_ext_flash_s1;
  input            cpu_instruction_master_granted_onchip_memory_s1;
  input            cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_instruction_master_qualified_request_descriptor_memory_s1;
  input            cpu_instruction_master_qualified_request_ext_flash_s1;
  input            cpu_instruction_master_qualified_request_onchip_memory_s1;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_instruction_master_read_data_valid_descriptor_memory_s1;
  input            cpu_instruction_master_read_data_valid_ext_flash_s1;
  input            cpu_instruction_master_read_data_valid_onchip_memory_s1;
  input            cpu_instruction_master_requests_cpu_jtag_debug_module;
  input            cpu_instruction_master_requests_descriptor_memory_s1;
  input            cpu_instruction_master_requests_ext_flash_s1;
  input            cpu_instruction_master_requests_onchip_memory_s1;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_descriptor_memory_s1_end_xfer;
  input            d1_flash_tristate_bridge_avalon_slave_end_xfer;
  input            d1_onchip_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            ext_flash_s1_wait_counter_eq_0;
  input   [ 15: 0] incoming_flash_tristate_bridge_data;
  input   [ 31: 0] onchip_memory_s1_readdata_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 30: 0] cpu_instruction_master_address_last_time;
  wire    [ 30: 0] cpu_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_instruction_master_dbs_address;
  wire    [  1: 0] cpu_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg     [  1: 0] cpu_instruction_master_latency_counter;
  wire    [  1: 0] cpu_instruction_master_next_dbs_rdv_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [  1: 0] p1_cpu_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_requests_cpu_jtag_debug_module) & (cpu_instruction_master_granted_cpu_jtag_debug_module | ~cpu_instruction_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_instruction_master_read))) & 1 & (cpu_instruction_master_qualified_request_descriptor_memory_s1 | ~cpu_instruction_master_requests_descriptor_memory_s1) & (cpu_instruction_master_granted_descriptor_memory_s1 | ~cpu_instruction_master_qualified_request_descriptor_memory_s1) & ((~cpu_instruction_master_qualified_request_descriptor_memory_s1 | ~(cpu_instruction_master_read) | (1 & (cpu_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_instruction_master_qualified_request_ext_flash_s1 | ~cpu_instruction_master_requests_ext_flash_s1) & (cpu_instruction_master_granted_ext_flash_s1 | ~cpu_instruction_master_qualified_request_ext_flash_s1) & ((~cpu_instruction_master_qualified_request_ext_flash_s1 | ~cpu_instruction_master_read | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & (cpu_instruction_master_dbs_address[1]) & cpu_instruction_master_read))) & 1 & (cpu_instruction_master_qualified_request_onchip_memory_s1 | ~cpu_instruction_master_requests_onchip_memory_s1) & (cpu_instruction_master_granted_onchip_memory_s1 | ~cpu_instruction_master_qualified_request_onchip_memory_s1) & ((~cpu_instruction_master_qualified_request_onchip_memory_s1 | ~(cpu_instruction_master_read) | (1 & (cpu_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = {3'b100,
    cpu_instruction_master_address[27 : 0]};

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_cpu_jtag_debug_module |
    cpu_instruction_master_granted_descriptor_memory_s1 |
    cpu_instruction_master_granted_ext_flash_s1 |
    cpu_instruction_master_granted_onchip_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_descriptor_memory_s1 |
    (cpu_instruction_master_read_data_valid_ext_flash_s1 & dbs_rdv_counter_overflow) |
    cpu_instruction_master_read_data_valid_onchip_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_data_valid_cpu_jtag_debug_module |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~(cpu_instruction_master_qualified_request_cpu_jtag_debug_module & cpu_instruction_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_descriptor_memory_s1}} | descriptor_memory_s1_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_ext_flash_s1}} | {incoming_flash_tristate_bridge_data[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~cpu_instruction_master_read_data_valid_onchip_memory_s1}} | onchip_memory_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {cpu_instruction_master_requests_descriptor_memory_s1}} & 1) |
    ({2 {cpu_instruction_master_requests_ext_flash_s1}} & 2) |
    ({2 {cpu_instruction_master_requests_onchip_memory_s1}} & 1);

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = incoming_flash_tristate_bridge_data;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_instruction_master_dbs_increment = (cpu_instruction_master_requests_ext_flash_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_instruction_master_dbs_address + cpu_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_instruction_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_instruction_master_next_dbs_rdv_counter = cpu_instruction_master_dbs_rdv_counter + cpu_instruction_master_dbs_rdv_counter_inc;

  //cpu_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_instruction_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_instruction_master_read_data_valid_ext_flash_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_instruction_master_dbs_rdv_counter <= cpu_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_instruction_master_dbs_rdv_counter[1] & ~cpu_instruction_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = cpu_instruction_master_granted_ext_flash_s1 & cpu_instruction_master_read & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer});


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_ddr2_s1_module (
                                            // inputs:
                                             clear_fifo,
                                             clk,
                                             data_in,
                                             read,
                                             reset_n,
                                             sync_reset,
                                             write,

                                            // outputs:
                                             data_out,
                                             empty,
                                             fifo_contains_ones_n,
                                             full
                                          )
;

  output  [  2: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  2: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  2: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  2: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  2: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  2: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  2: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  2: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  2: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  2: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  2: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  2: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  2: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  2: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  2: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  2: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  2: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  2: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  2: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  2: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  2: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  2: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  2: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  2: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  2: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  2: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  2: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  2: 0] p31_stage_31;
  wire             p3_full_3;
  wire    [  2: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  2: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  2: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  2: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  2: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  2: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  2: 0] p9_stage_9;
  reg     [  2: 0] stage_0;
  reg     [  2: 0] stage_1;
  reg     [  2: 0] stage_10;
  reg     [  2: 0] stage_11;
  reg     [  2: 0] stage_12;
  reg     [  2: 0] stage_13;
  reg     [  2: 0] stage_14;
  reg     [  2: 0] stage_15;
  reg     [  2: 0] stage_16;
  reg     [  2: 0] stage_17;
  reg     [  2: 0] stage_18;
  reg     [  2: 0] stage_19;
  reg     [  2: 0] stage_2;
  reg     [  2: 0] stage_20;
  reg     [  2: 0] stage_21;
  reg     [  2: 0] stage_22;
  reg     [  2: 0] stage_23;
  reg     [  2: 0] stage_24;
  reg     [  2: 0] stage_25;
  reg     [  2: 0] stage_26;
  reg     [  2: 0] stage_27;
  reg     [  2: 0] stage_28;
  reg     [  2: 0] stage_29;
  reg     [  2: 0] stage_3;
  reg     [  2: 0] stage_30;
  reg     [  2: 0] stage_31;
  reg     [  2: 0] stage_4;
  reg     [  2: 0] stage_5;
  reg     [  2: 0] stage_6;
  reg     [  2: 0] stage_7;
  reg     [  2: 0] stage_8;
  reg     [  2: 0] stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_SS_OCT_SOPC_burst_0_downstream_to_ddr2_s1_module (
                                                                       // inputs:
                                                                        clear_fifo,
                                                                        clk,
                                                                        data_in,
                                                                        read,
                                                                        reset_n,
                                                                        sync_reset,
                                                                        write,

                                                                       // outputs:
                                                                        data_out,
                                                                        empty,
                                                                        fifo_contains_ones_n,
                                                                        full
                                                                     )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pipeline_bridge_ddr2_m1_to_ddr2_s1_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr2_s1_arbitrator (
                            // inputs:
                             SS_OCT_SOPC_burst_0_downstream_address_to_slave,
                             SS_OCT_SOPC_burst_0_downstream_arbitrationshare,
                             SS_OCT_SOPC_burst_0_downstream_burstcount,
                             SS_OCT_SOPC_burst_0_downstream_byteenable,
                             SS_OCT_SOPC_burst_0_downstream_latency_counter,
                             SS_OCT_SOPC_burst_0_downstream_read,
                             SS_OCT_SOPC_burst_0_downstream_write,
                             SS_OCT_SOPC_burst_0_downstream_writedata,
                             clk,
                             ddr2_s1_readdata,
                             ddr2_s1_readdatavalid,
                             ddr2_s1_resetrequest_n,
                             ddr2_s1_waitrequest_n,
                             pipeline_bridge_ddr2_m1_address_to_slave,
                             pipeline_bridge_ddr2_m1_burstcount,
                             pipeline_bridge_ddr2_m1_byteenable,
                             pipeline_bridge_ddr2_m1_chipselect,
                             pipeline_bridge_ddr2_m1_latency_counter,
                             pipeline_bridge_ddr2_m1_read,
                             pipeline_bridge_ddr2_m1_write,
                             pipeline_bridge_ddr2_m1_writedata,
                             reset_n,

                            // outputs:
                             SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1,
                             SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1,
                             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1,
                             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register,
                             SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1,
                             d1_ddr2_s1_end_xfer,
                             ddr2_s1_address,
                             ddr2_s1_beginbursttransfer,
                             ddr2_s1_burstcount,
                             ddr2_s1_byteenable,
                             ddr2_s1_read,
                             ddr2_s1_readdata_from_sa,
                             ddr2_s1_resetrequest_n_from_sa,
                             ddr2_s1_waitrequest_n_from_sa,
                             ddr2_s1_write,
                             ddr2_s1_writedata,
                             pipeline_bridge_ddr2_m1_granted_ddr2_s1,
                             pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1,
                             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1,
                             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register,
                             pipeline_bridge_ddr2_m1_requests_ddr2_s1
                          )
;

  output           SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1;
  output           SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1;
  output           SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1;
  output           SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register;
  output           SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1;
  output           d1_ddr2_s1_end_xfer;
  output  [ 24: 0] ddr2_s1_address;
  output           ddr2_s1_beginbursttransfer;
  output  [  2: 0] ddr2_s1_burstcount;
  output  [ 31: 0] ddr2_s1_byteenable;
  output           ddr2_s1_read;
  output  [255: 0] ddr2_s1_readdata_from_sa;
  output           ddr2_s1_resetrequest_n_from_sa;
  output           ddr2_s1_waitrequest_n_from_sa;
  output           ddr2_s1_write;
  output  [255: 0] ddr2_s1_writedata;
  output           pipeline_bridge_ddr2_m1_granted_ddr2_s1;
  output           pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1;
  output           pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;
  output           pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register;
  output           pipeline_bridge_ddr2_m1_requests_ddr2_s1;
  input   [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address_to_slave;
  input   [  3: 0] SS_OCT_SOPC_burst_0_downstream_arbitrationshare;
  input   [  2: 0] SS_OCT_SOPC_burst_0_downstream_burstcount;
  input   [ 31: 0] SS_OCT_SOPC_burst_0_downstream_byteenable;
  input            SS_OCT_SOPC_burst_0_downstream_latency_counter;
  input            SS_OCT_SOPC_burst_0_downstream_read;
  input            SS_OCT_SOPC_burst_0_downstream_write;
  input   [255: 0] SS_OCT_SOPC_burst_0_downstream_writedata;
  input            clk;
  input   [255: 0] ddr2_s1_readdata;
  input            ddr2_s1_readdatavalid;
  input            ddr2_s1_resetrequest_n;
  input            ddr2_s1_waitrequest_n;
  input   [ 29: 0] pipeline_bridge_ddr2_m1_address_to_slave;
  input            pipeline_bridge_ddr2_m1_burstcount;
  input   [  3: 0] pipeline_bridge_ddr2_m1_byteenable;
  input            pipeline_bridge_ddr2_m1_chipselect;
  input            pipeline_bridge_ddr2_m1_latency_counter;
  input            pipeline_bridge_ddr2_m1_read;
  input            pipeline_bridge_ddr2_m1_write;
  input   [ 31: 0] pipeline_bridge_ddr2_m1_writedata;
  input            reset_n;

  wire             SS_OCT_SOPC_burst_0_downstream_arbiterlock;
  wire             SS_OCT_SOPC_burst_0_downstream_arbiterlock2;
  wire             SS_OCT_SOPC_burst_0_downstream_continuerequest;
  wire             SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_rdv_fifo_empty_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_rdv_fifo_output_from_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register;
  wire             SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1;
  reg              d1_ddr2_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 24: 0] ddr2_s1_address;
  wire             ddr2_s1_allgrants;
  wire             ddr2_s1_allow_new_arb_cycle;
  wire             ddr2_s1_any_bursting_master_saved_grant;
  wire             ddr2_s1_any_continuerequest;
  reg     [  1: 0] ddr2_s1_arb_addend;
  wire             ddr2_s1_arb_counter_enable;
  reg     [  3: 0] ddr2_s1_arb_share_counter;
  wire    [  3: 0] ddr2_s1_arb_share_counter_next_value;
  wire    [  3: 0] ddr2_s1_arb_share_set_values;
  wire    [  1: 0] ddr2_s1_arb_winner;
  wire             ddr2_s1_arbitration_holdoff_internal;
  reg     [  1: 0] ddr2_s1_bbt_burstcounter;
  wire             ddr2_s1_beginbursttransfer;
  wire             ddr2_s1_beginbursttransfer_internal;
  wire             ddr2_s1_begins_xfer;
  wire    [  2: 0] ddr2_s1_burstcount;
  wire             ddr2_s1_burstcount_fifo_empty;
  wire    [ 31: 0] ddr2_s1_byteenable;
  wire    [  3: 0] ddr2_s1_chosen_master_double_vector;
  wire    [  1: 0] ddr2_s1_chosen_master_rot_left;
  reg     [  2: 0] ddr2_s1_current_burst;
  wire    [  2: 0] ddr2_s1_current_burst_minus_one;
  wire             ddr2_s1_end_xfer;
  wire             ddr2_s1_firsttransfer;
  wire    [  1: 0] ddr2_s1_grant_vector;
  wire             ddr2_s1_in_a_read_cycle;
  wire             ddr2_s1_in_a_write_cycle;
  reg              ddr2_s1_load_fifo;
  wire    [  1: 0] ddr2_s1_master_qreq_vector;
  wire             ddr2_s1_move_on_to_next_transaction;
  wire    [  1: 0] ddr2_s1_next_bbt_burstcount;
  wire    [  2: 0] ddr2_s1_next_burst_count;
  wire             ddr2_s1_non_bursting_master_requests;
  wire             ddr2_s1_read;
  wire    [255: 0] ddr2_s1_readdata_from_sa;
  wire             ddr2_s1_readdatavalid_from_sa;
  reg              ddr2_s1_reg_firsttransfer;
  wire             ddr2_s1_resetrequest_n_from_sa;
  reg     [  1: 0] ddr2_s1_saved_chosen_master_vector;
  wire    [  2: 0] ddr2_s1_selected_burstcount;
  reg              ddr2_s1_slavearbiterlockenable;
  wire             ddr2_s1_slavearbiterlockenable2;
  wire             ddr2_s1_this_cycle_is_the_last_burst;
  wire    [  2: 0] ddr2_s1_transaction_burst_count;
  wire             ddr2_s1_unreg_firsttransfer;
  wire             ddr2_s1_waitrequest_n_from_sa;
  wire             ddr2_s1_waits_for_read;
  wire             ddr2_s1_waits_for_write;
  wire             ddr2_s1_write;
  wire    [255: 0] ddr2_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ddr2_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_SS_OCT_SOPC_burst_0_downstream_granted_slave_ddr2_s1;
  reg              last_cycle_pipeline_bridge_ddr2_m1_granted_slave_ddr2_s1;
  wire             p0_ddr2_s1_load_fifo;
  wire             pipeline_bridge_ddr2_m1_arbiterlock;
  wire             pipeline_bridge_ddr2_m1_arbiterlock2;
  wire    [ 31: 0] pipeline_bridge_ddr2_m1_byteenable_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_continuerequest;
  wire             pipeline_bridge_ddr2_m1_granted_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_rdv_fifo_empty_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_rdv_fifo_output_from_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register;
  wire             pipeline_bridge_ddr2_m1_requests_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_saved_grant_ddr2_s1;
  wire    [255: 0] pipeline_bridge_ddr2_m1_writedata_replicated;
  wire    [ 29: 0] shifted_address_to_ddr2_s1_from_SS_OCT_SOPC_burst_0_downstream;
  wire    [ 29: 0] shifted_address_to_ddr2_s1_from_pipeline_bridge_ddr2_m1;
  wire             wait_for_ddr2_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ddr2_s1_end_xfer;
    end


  assign ddr2_s1_begins_xfer = ~d1_reasons_to_wait & ((SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1 | pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1));
  //assign ddr2_s1_readdata_from_sa = ddr2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_s1_readdata_from_sa = ddr2_s1_readdata;

  assign SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1 = (1) & (SS_OCT_SOPC_burst_0_downstream_read | SS_OCT_SOPC_burst_0_downstream_write);
  //assign ddr2_s1_waitrequest_n_from_sa = ddr2_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_s1_waitrequest_n_from_sa = ddr2_s1_waitrequest_n;

  //assign ddr2_s1_readdatavalid_from_sa = ddr2_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_s1_readdatavalid_from_sa = ddr2_s1_readdatavalid;

  //ddr2_s1_arb_share_counter set values, which is an e_mux
  assign ddr2_s1_arb_share_set_values = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_arbitrationshare :
    (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_arbitrationshare :
    1;

  //ddr2_s1_non_bursting_master_requests mux, which is an e_mux
  assign ddr2_s1_non_bursting_master_requests = 0 |
    pipeline_bridge_ddr2_m1_requests_ddr2_s1 |
    pipeline_bridge_ddr2_m1_requests_ddr2_s1;

  //ddr2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ddr2_s1_any_bursting_master_saved_grant = SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1 |
    SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1;

  //ddr2_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ddr2_s1_arb_share_counter_next_value = ddr2_s1_firsttransfer ? (ddr2_s1_arb_share_set_values - 1) : |ddr2_s1_arb_share_counter ? (ddr2_s1_arb_share_counter - 1) : 0;

  //ddr2_s1_allgrants all slave grants, which is an e_mux
  assign ddr2_s1_allgrants = (|ddr2_s1_grant_vector) |
    (|ddr2_s1_grant_vector) |
    (|ddr2_s1_grant_vector) |
    (|ddr2_s1_grant_vector);

  //ddr2_s1_end_xfer assignment, which is an e_assign
  assign ddr2_s1_end_xfer = ~(ddr2_s1_waits_for_read | ddr2_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ddr2_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ddr2_s1 = ddr2_s1_end_xfer & (~ddr2_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ddr2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ddr2_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ddr2_s1 & ddr2_s1_allgrants) | (end_xfer_arb_share_counter_term_ddr2_s1 & ~ddr2_s1_non_bursting_master_requests);

  //ddr2_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_arb_share_counter <= 0;
      else if (ddr2_s1_arb_counter_enable)
          ddr2_s1_arb_share_counter <= ddr2_s1_arb_share_counter_next_value;
    end


  //ddr2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_slavearbiterlockenable <= 0;
      else if ((|ddr2_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ddr2_s1) | (end_xfer_arb_share_counter_term_ddr2_s1 & ~ddr2_s1_non_bursting_master_requests))
          ddr2_s1_slavearbiterlockenable <= |ddr2_s1_arb_share_counter_next_value;
    end


  //SS_OCT_SOPC_burst_0/downstream ddr2/s1 arbiterlock, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_arbiterlock = ddr2_s1_slavearbiterlockenable & SS_OCT_SOPC_burst_0_downstream_continuerequest;

  //ddr2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ddr2_s1_slavearbiterlockenable2 = |ddr2_s1_arb_share_counter_next_value;

  //SS_OCT_SOPC_burst_0/downstream ddr2/s1 arbiterlock2, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_arbiterlock2 = ddr2_s1_slavearbiterlockenable2 & SS_OCT_SOPC_burst_0_downstream_continuerequest;

  //pipeline_bridge_ddr2/m1 ddr2/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_ddr2_m1_arbiterlock = ddr2_s1_slavearbiterlockenable & pipeline_bridge_ddr2_m1_continuerequest;

  //pipeline_bridge_ddr2/m1 ddr2/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_ddr2_m1_arbiterlock2 = ddr2_s1_slavearbiterlockenable2 & pipeline_bridge_ddr2_m1_continuerequest;

  //pipeline_bridge_ddr2/m1 granted ddr2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pipeline_bridge_ddr2_m1_granted_slave_ddr2_s1 <= 0;
      else 
        last_cycle_pipeline_bridge_ddr2_m1_granted_slave_ddr2_s1 <= pipeline_bridge_ddr2_m1_saved_grant_ddr2_s1 ? 1 : (ddr2_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_pipeline_bridge_ddr2_m1_granted_slave_ddr2_s1;
    end


  //pipeline_bridge_ddr2_m1_continuerequest continued request, which is an e_mux
  assign pipeline_bridge_ddr2_m1_continuerequest = last_cycle_pipeline_bridge_ddr2_m1_granted_slave_ddr2_s1 & pipeline_bridge_ddr2_m1_requests_ddr2_s1;

  //ddr2_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ddr2_s1_any_continuerequest = pipeline_bridge_ddr2_m1_continuerequest |
    SS_OCT_SOPC_burst_0_downstream_continuerequest;

  assign SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1 = SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1 & ~((SS_OCT_SOPC_burst_0_downstream_read & ((SS_OCT_SOPC_burst_0_downstream_latency_counter != 0) | (1 < SS_OCT_SOPC_burst_0_downstream_latency_counter))) | pipeline_bridge_ddr2_m1_arbiterlock);
  //unique name for ddr2_s1_move_on_to_next_transaction, which is an e_assign
  assign ddr2_s1_move_on_to_next_transaction = ddr2_s1_this_cycle_is_the_last_burst & ddr2_s1_load_fifo;

  //the currently selected burstcount for ddr2_s1, which is an e_mux
  assign ddr2_s1_selected_burstcount = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_burstcount :
    1;

  //burstcount_fifo_for_ddr2_s1, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_ddr2_s1_module burstcount_fifo_for_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (ddr2_s1_selected_burstcount),
      .data_out             (ddr2_s1_transaction_burst_count),
      .empty                (ddr2_s1_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (ddr2_s1_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr2_s1_waits_for_read & ddr2_s1_load_fifo & ~(ddr2_s1_this_cycle_is_the_last_burst & ddr2_s1_burstcount_fifo_empty))
    );

  //ddr2_s1 current burst minus one, which is an e_assign
  assign ddr2_s1_current_burst_minus_one = ddr2_s1_current_burst - 1;

  //what to load in current_burst, for ddr2_s1, which is an e_mux
  assign ddr2_s1_next_burst_count = (((in_a_read_cycle & ~ddr2_s1_waits_for_read) & ~ddr2_s1_load_fifo))? ddr2_s1_selected_burstcount :
    ((in_a_read_cycle & ~ddr2_s1_waits_for_read & ddr2_s1_this_cycle_is_the_last_burst & ddr2_s1_burstcount_fifo_empty))? ddr2_s1_selected_burstcount :
    (ddr2_s1_this_cycle_is_the_last_burst)? ddr2_s1_transaction_burst_count :
    ddr2_s1_current_burst_minus_one;

  //the current burst count for ddr2_s1, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_current_burst <= 0;
      else if (ddr2_s1_readdatavalid_from_sa | (~ddr2_s1_load_fifo & (in_a_read_cycle & ~ddr2_s1_waits_for_read)))
          ddr2_s1_current_burst <= ddr2_s1_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_ddr2_s1_load_fifo = (~ddr2_s1_load_fifo)? 1 :
    (((in_a_read_cycle & ~ddr2_s1_waits_for_read) & ddr2_s1_load_fifo))? 1 :
    ~ddr2_s1_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_load_fifo <= 0;
      else if ((in_a_read_cycle & ~ddr2_s1_waits_for_read) & ~ddr2_s1_load_fifo | ddr2_s1_this_cycle_is_the_last_burst)
          ddr2_s1_load_fifo <= p0_ddr2_s1_load_fifo;
    end


  //the last cycle in the burst for ddr2_s1, which is an e_assign
  assign ddr2_s1_this_cycle_is_the_last_burst = ~(|ddr2_s1_current_burst_minus_one) & ddr2_s1_readdatavalid_from_sa;

  //rdv_fifo_for_SS_OCT_SOPC_burst_0_downstream_to_ddr2_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_SS_OCT_SOPC_burst_0_downstream_to_ddr2_s1_module rdv_fifo_for_SS_OCT_SOPC_burst_0_downstream_to_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1),
      .data_out             (SS_OCT_SOPC_burst_0_downstream_rdv_fifo_output_from_ddr2_s1),
      .empty                (),
      .fifo_contains_ones_n (SS_OCT_SOPC_burst_0_downstream_rdv_fifo_empty_ddr2_s1),
      .full                 (),
      .read                 (ddr2_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr2_s1_waits_for_read)
    );

  assign SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register = ~SS_OCT_SOPC_burst_0_downstream_rdv_fifo_empty_ddr2_s1;
  //local readdatavalid SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1, which is an e_mux
  assign SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1 = (ddr2_s1_readdatavalid_from_sa & SS_OCT_SOPC_burst_0_downstream_rdv_fifo_output_from_ddr2_s1) & ~ SS_OCT_SOPC_burst_0_downstream_rdv_fifo_empty_ddr2_s1;

  //ddr2_s1_writedata mux, which is an e_mux
  assign ddr2_s1_writedata = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_writedata :
    pipeline_bridge_ddr2_m1_writedata_replicated;

  assign pipeline_bridge_ddr2_m1_requests_ddr2_s1 = (1) & pipeline_bridge_ddr2_m1_chipselect;
  //SS_OCT_SOPC_burst_0/downstream granted ddr2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_SS_OCT_SOPC_burst_0_downstream_granted_slave_ddr2_s1 <= 0;
      else 
        last_cycle_SS_OCT_SOPC_burst_0_downstream_granted_slave_ddr2_s1 <= SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1 ? 1 : (ddr2_s1_arbitration_holdoff_internal | ~SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1) ? 0 : last_cycle_SS_OCT_SOPC_burst_0_downstream_granted_slave_ddr2_s1;
    end


  //SS_OCT_SOPC_burst_0_downstream_continuerequest continued request, which is an e_mux
  assign SS_OCT_SOPC_burst_0_downstream_continuerequest = last_cycle_SS_OCT_SOPC_burst_0_downstream_granted_slave_ddr2_s1 & 1;

  assign pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1 = pipeline_bridge_ddr2_m1_requests_ddr2_s1 & ~(((pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect) & ((pipeline_bridge_ddr2_m1_latency_counter != 0) | (1 < pipeline_bridge_ddr2_m1_latency_counter))) | SS_OCT_SOPC_burst_0_downstream_arbiterlock);
  //rdv_fifo_for_pipeline_bridge_ddr2_m1_to_ddr2_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pipeline_bridge_ddr2_m1_to_ddr2_s1_module rdv_fifo_for_pipeline_bridge_ddr2_m1_to_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_ddr2_m1_granted_ddr2_s1),
      .data_out             (pipeline_bridge_ddr2_m1_rdv_fifo_output_from_ddr2_s1),
      .empty                (),
      .fifo_contains_ones_n (pipeline_bridge_ddr2_m1_rdv_fifo_empty_ddr2_s1),
      .full                 (),
      .read                 (ddr2_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr2_s1_waits_for_read)
    );

  assign pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register = ~pipeline_bridge_ddr2_m1_rdv_fifo_empty_ddr2_s1;
  //local readdatavalid pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1, which is an e_mux
  assign pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1 = (ddr2_s1_readdatavalid_from_sa & pipeline_bridge_ddr2_m1_rdv_fifo_output_from_ddr2_s1) & ~ pipeline_bridge_ddr2_m1_rdv_fifo_empty_ddr2_s1;

  //replicate narrow data for wide slave
  assign pipeline_bridge_ddr2_m1_writedata_replicated = {pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata,
    pipeline_bridge_ddr2_m1_writedata};

  //allow new arb cycle for ddr2/s1, which is an e_assign
  assign ddr2_s1_allow_new_arb_cycle = ~SS_OCT_SOPC_burst_0_downstream_arbiterlock & ~pipeline_bridge_ddr2_m1_arbiterlock;

  //pipeline_bridge_ddr2/m1 assignment into master qualified-requests vector for ddr2/s1, which is an e_assign
  assign ddr2_s1_master_qreq_vector[0] = pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1;

  //pipeline_bridge_ddr2/m1 grant ddr2/s1, which is an e_assign
  assign pipeline_bridge_ddr2_m1_granted_ddr2_s1 = ddr2_s1_grant_vector[0];

  //pipeline_bridge_ddr2/m1 saved-grant ddr2/s1, which is an e_assign
  assign pipeline_bridge_ddr2_m1_saved_grant_ddr2_s1 = ddr2_s1_arb_winner[0] && pipeline_bridge_ddr2_m1_requests_ddr2_s1;

  //SS_OCT_SOPC_burst_0/downstream assignment into master qualified-requests vector for ddr2/s1, which is an e_assign
  assign ddr2_s1_master_qreq_vector[1] = SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1;

  //SS_OCT_SOPC_burst_0/downstream grant ddr2/s1, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 = ddr2_s1_grant_vector[1];

  //SS_OCT_SOPC_burst_0/downstream saved-grant ddr2/s1, which is an e_assign
  assign SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1 = ddr2_s1_arb_winner[1];

  //ddr2/s1 chosen-master double-vector, which is an e_assign
  assign ddr2_s1_chosen_master_double_vector = {ddr2_s1_master_qreq_vector, ddr2_s1_master_qreq_vector} & ({~ddr2_s1_master_qreq_vector, ~ddr2_s1_master_qreq_vector} + ddr2_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign ddr2_s1_arb_winner = (ddr2_s1_allow_new_arb_cycle & | ddr2_s1_grant_vector) ? ddr2_s1_grant_vector : ddr2_s1_saved_chosen_master_vector;

  //saved ddr2_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_saved_chosen_master_vector <= 0;
      else if (ddr2_s1_allow_new_arb_cycle)
          ddr2_s1_saved_chosen_master_vector <= |ddr2_s1_grant_vector ? ddr2_s1_grant_vector : ddr2_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ddr2_s1_grant_vector = {(ddr2_s1_chosen_master_double_vector[1] | ddr2_s1_chosen_master_double_vector[3]),
    (ddr2_s1_chosen_master_double_vector[0] | ddr2_s1_chosen_master_double_vector[2])};

  //ddr2/s1 chosen master rotated left, which is an e_assign
  assign ddr2_s1_chosen_master_rot_left = (ddr2_s1_arb_winner << 1) ? (ddr2_s1_arb_winner << 1) : 1;

  //ddr2/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_arb_addend <= 1;
      else if (|ddr2_s1_grant_vector)
          ddr2_s1_arb_addend <= ddr2_s1_end_xfer? ddr2_s1_chosen_master_rot_left : ddr2_s1_grant_vector;
    end


  //assign ddr2_s1_resetrequest_n_from_sa = ddr2_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_s1_resetrequest_n_from_sa = ddr2_s1_resetrequest_n;

  //ddr2_s1_firsttransfer first transaction, which is an e_assign
  assign ddr2_s1_firsttransfer = ddr2_s1_begins_xfer ? ddr2_s1_unreg_firsttransfer : ddr2_s1_reg_firsttransfer;

  //ddr2_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ddr2_s1_unreg_firsttransfer = ~(ddr2_s1_slavearbiterlockenable & ddr2_s1_any_continuerequest);

  //ddr2_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_reg_firsttransfer <= 1'b1;
      else if (ddr2_s1_begins_xfer)
          ddr2_s1_reg_firsttransfer <= ddr2_s1_unreg_firsttransfer;
    end


  //ddr2_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign ddr2_s1_next_bbt_burstcount = ((((ddr2_s1_write) && (ddr2_s1_bbt_burstcounter == 0))))? (ddr2_s1_burstcount - 1) :
    ((((ddr2_s1_read) && (ddr2_s1_bbt_burstcounter == 0))))? 0 :
    (ddr2_s1_bbt_burstcounter - 1);

  //ddr2_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_s1_bbt_burstcounter <= 0;
      else if (ddr2_s1_begins_xfer)
          ddr2_s1_bbt_burstcounter <= ddr2_s1_next_bbt_burstcount;
    end


  //ddr2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ddr2_s1_beginbursttransfer_internal = ddr2_s1_begins_xfer & (ddr2_s1_bbt_burstcounter == 0);

  //ddr2/s1 begin burst transfer to slave, which is an e_assign
  assign ddr2_s1_beginbursttransfer = ddr2_s1_beginbursttransfer_internal;

  //ddr2_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ddr2_s1_arbitration_holdoff_internal = ddr2_s1_begins_xfer & ddr2_s1_firsttransfer;

  //ddr2_s1_read assignment, which is an e_mux
  assign ddr2_s1_read = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 & SS_OCT_SOPC_burst_0_downstream_read) | (pipeline_bridge_ddr2_m1_granted_ddr2_s1 & (pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect));

  //ddr2_s1_write assignment, which is an e_mux
  assign ddr2_s1_write = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 & SS_OCT_SOPC_burst_0_downstream_write) | (pipeline_bridge_ddr2_m1_granted_ddr2_s1 & (pipeline_bridge_ddr2_m1_write & pipeline_bridge_ddr2_m1_chipselect));

  assign shifted_address_to_ddr2_s1_from_SS_OCT_SOPC_burst_0_downstream = SS_OCT_SOPC_burst_0_downstream_address_to_slave;
  //ddr2_s1_address mux, which is an e_mux
  assign ddr2_s1_address = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? (shifted_address_to_ddr2_s1_from_SS_OCT_SOPC_burst_0_downstream >> 5) :
    (shifted_address_to_ddr2_s1_from_pipeline_bridge_ddr2_m1 >> 5);

  assign shifted_address_to_ddr2_s1_from_pipeline_bridge_ddr2_m1 = pipeline_bridge_ddr2_m1_address_to_slave;
  //d1_ddr2_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ddr2_s1_end_xfer <= 1;
      else 
        d1_ddr2_s1_end_xfer <= ddr2_s1_end_xfer;
    end


  //ddr2_s1_waits_for_read in a cycle, which is an e_mux
  assign ddr2_s1_waits_for_read = ddr2_s1_in_a_read_cycle & ~ddr2_s1_waitrequest_n_from_sa;

  //ddr2_s1_in_a_read_cycle assignment, which is an e_assign
  assign ddr2_s1_in_a_read_cycle = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 & SS_OCT_SOPC_burst_0_downstream_read) | (pipeline_bridge_ddr2_m1_granted_ddr2_s1 & (pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect));

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ddr2_s1_in_a_read_cycle;

  //ddr2_s1_waits_for_write in a cycle, which is an e_mux
  assign ddr2_s1_waits_for_write = ddr2_s1_in_a_write_cycle & ~ddr2_s1_waitrequest_n_from_sa;

  //ddr2_s1_in_a_write_cycle assignment, which is an e_assign
  assign ddr2_s1_in_a_write_cycle = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 & SS_OCT_SOPC_burst_0_downstream_write) | (pipeline_bridge_ddr2_m1_granted_ddr2_s1 & (pipeline_bridge_ddr2_m1_write & pipeline_bridge_ddr2_m1_chipselect));

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ddr2_s1_in_a_write_cycle;

  assign wait_for_ddr2_s1_counter = 0;
  //ddr2_s1_byteenable byte enable port mux, which is an e_mux
  assign ddr2_s1_byteenable = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_byteenable :
    (pipeline_bridge_ddr2_m1_granted_ddr2_s1)? pipeline_bridge_ddr2_m1_byteenable_ddr2_s1 :
    -1;

  //byte_enable_mux for pipeline_bridge_ddr2/m1 and ddr2/s1, which is an e_mux
  assign pipeline_bridge_ddr2_m1_byteenable_ddr2_s1 = (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 0)? pipeline_bridge_ddr2_m1_byteenable :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 1)? {pipeline_bridge_ddr2_m1_byteenable, {4'b0}} :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 2)? {pipeline_bridge_ddr2_m1_byteenable, {8'b0}} :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 3)? {pipeline_bridge_ddr2_m1_byteenable, {12'b0}} :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 4)? {pipeline_bridge_ddr2_m1_byteenable, {16'b0}} :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 5)? {pipeline_bridge_ddr2_m1_byteenable, {20'b0}} :
    (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2] == 6)? {pipeline_bridge_ddr2_m1_byteenable, {24'b0}} :
    {pipeline_bridge_ddr2_m1_byteenable, {28'b0}};

  //burstcount mux, which is an e_mux
  assign ddr2_s1_burstcount = (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1)? SS_OCT_SOPC_burst_0_downstream_burstcount :
    (pipeline_bridge_ddr2_m1_granted_ddr2_s1)? pipeline_bridge_ddr2_m1_burstcount :
    1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //SS_OCT_SOPC_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1 && (SS_OCT_SOPC_burst_0_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave ddr2/s1", $time);
          $stop;
        end
    end


  //SS_OCT_SOPC_burst_0/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1 && (SS_OCT_SOPC_burst_0_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: SS_OCT_SOPC_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave ddr2/s1", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_ddr2_m1_requests_ddr2_s1 && (pipeline_bridge_ddr2_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge_ddr2/m1 drove 0 on its 'burstcount' port while accessing slave ddr2/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1 + pipeline_bridge_ddr2_m1_granted_ddr2_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (SS_OCT_SOPC_burst_0_downstream_saved_grant_ddr2_s1 + pipeline_bridge_ddr2_m1_saved_grant_ddr2_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_reset_clk_50_domain_synch_module (
                                                      // inputs:
                                                       clk,
                                                       data_in,
                                                       reset_n,

                                                      // outputs:
                                                       data_out
                                                    )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module descriptor_memory_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          cpu_data_master_address_to_slave,
                                          cpu_data_master_byteenable,
                                          cpu_data_master_latency_counter,
                                          cpu_data_master_read,
                                          cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                          cpu_data_master_write,
                                          cpu_data_master_writedata,
                                          cpu_instruction_master_address_to_slave,
                                          cpu_instruction_master_latency_counter,
                                          cpu_instruction_master_read,
                                          descriptor_memory_s1_readdata,
                                          reset_n,
                                          sgdma_rx_descriptor_read_address_to_slave,
                                          sgdma_rx_descriptor_read_latency_counter,
                                          sgdma_rx_descriptor_read_read,
                                          sgdma_rx_descriptor_write_address_to_slave,
                                          sgdma_rx_descriptor_write_write,
                                          sgdma_rx_descriptor_write_writedata,
                                          sgdma_tx_descriptor_read_address_to_slave,
                                          sgdma_tx_descriptor_read_latency_counter,
                                          sgdma_tx_descriptor_read_read,
                                          sgdma_tx_descriptor_write_address_to_slave,
                                          sgdma_tx_descriptor_write_write,
                                          sgdma_tx_descriptor_write_writedata,

                                         // outputs:
                                          cpu_data_master_granted_descriptor_memory_s1,
                                          cpu_data_master_qualified_request_descriptor_memory_s1,
                                          cpu_data_master_read_data_valid_descriptor_memory_s1,
                                          cpu_data_master_requests_descriptor_memory_s1,
                                          cpu_instruction_master_granted_descriptor_memory_s1,
                                          cpu_instruction_master_qualified_request_descriptor_memory_s1,
                                          cpu_instruction_master_read_data_valid_descriptor_memory_s1,
                                          cpu_instruction_master_requests_descriptor_memory_s1,
                                          d1_descriptor_memory_s1_end_xfer,
                                          descriptor_memory_s1_address,
                                          descriptor_memory_s1_byteenable,
                                          descriptor_memory_s1_chipselect,
                                          descriptor_memory_s1_clken,
                                          descriptor_memory_s1_readdata_from_sa,
                                          descriptor_memory_s1_write,
                                          descriptor_memory_s1_writedata,
                                          sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_requests_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_requests_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_requests_descriptor_memory_s1
                                       )
;

  output           cpu_data_master_granted_descriptor_memory_s1;
  output           cpu_data_master_qualified_request_descriptor_memory_s1;
  output           cpu_data_master_read_data_valid_descriptor_memory_s1;
  output           cpu_data_master_requests_descriptor_memory_s1;
  output           cpu_instruction_master_granted_descriptor_memory_s1;
  output           cpu_instruction_master_qualified_request_descriptor_memory_s1;
  output           cpu_instruction_master_read_data_valid_descriptor_memory_s1;
  output           cpu_instruction_master_requests_descriptor_memory_s1;
  output           d1_descriptor_memory_s1_end_xfer;
  output  [  8: 0] descriptor_memory_s1_address;
  output  [  3: 0] descriptor_memory_s1_byteenable;
  output           descriptor_memory_s1_chipselect;
  output           descriptor_memory_s1_clken;
  output  [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  output           descriptor_memory_s1_write;
  output  [ 31: 0] descriptor_memory_s1_writedata;
  output           sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 30: 0] cpu_instruction_master_address_to_slave;
  input   [  1: 0] cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input   [ 31: 0] descriptor_memory_s1_readdata;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  input            sgdma_rx_descriptor_read_latency_counter;
  input            sgdma_rx_descriptor_read_read;
  input   [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;
  input   [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  input            sgdma_tx_descriptor_read_latency_counter;
  input            sgdma_tx_descriptor_read_read;
  input   [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_descriptor_memory_s1;
  wire             cpu_data_master_qualified_request_descriptor_memory_s1;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1;
  reg              cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             cpu_data_master_requests_descriptor_memory_s1;
  wire             cpu_data_master_saved_grant_descriptor_memory_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_descriptor_memory_s1;
  wire             cpu_instruction_master_qualified_request_descriptor_memory_s1;
  wire             cpu_instruction_master_read_data_valid_descriptor_memory_s1;
  reg              cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             cpu_instruction_master_requests_descriptor_memory_s1;
  wire             cpu_instruction_master_saved_grant_descriptor_memory_s1;
  reg              d1_descriptor_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [  8: 0] descriptor_memory_s1_address;
  wire             descriptor_memory_s1_allgrants;
  wire             descriptor_memory_s1_allow_new_arb_cycle;
  wire             descriptor_memory_s1_any_bursting_master_saved_grant;
  wire             descriptor_memory_s1_any_continuerequest;
  reg     [  5: 0] descriptor_memory_s1_arb_addend;
  wire             descriptor_memory_s1_arb_counter_enable;
  reg     [  1: 0] descriptor_memory_s1_arb_share_counter;
  wire    [  1: 0] descriptor_memory_s1_arb_share_counter_next_value;
  wire    [  1: 0] descriptor_memory_s1_arb_share_set_values;
  wire    [  5: 0] descriptor_memory_s1_arb_winner;
  wire             descriptor_memory_s1_arbitration_holdoff_internal;
  wire             descriptor_memory_s1_beginbursttransfer_internal;
  wire             descriptor_memory_s1_begins_xfer;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire    [ 11: 0] descriptor_memory_s1_chosen_master_double_vector;
  wire    [  5: 0] descriptor_memory_s1_chosen_master_rot_left;
  wire             descriptor_memory_s1_clken;
  wire             descriptor_memory_s1_end_xfer;
  wire             descriptor_memory_s1_firsttransfer;
  wire    [  5: 0] descriptor_memory_s1_grant_vector;
  wire             descriptor_memory_s1_in_a_read_cycle;
  wire             descriptor_memory_s1_in_a_write_cycle;
  wire    [  5: 0] descriptor_memory_s1_master_qreq_vector;
  wire             descriptor_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  reg              descriptor_memory_s1_reg_firsttransfer;
  reg     [  5: 0] descriptor_memory_s1_saved_chosen_master_vector;
  reg              descriptor_memory_s1_slavearbiterlockenable;
  wire             descriptor_memory_s1_slavearbiterlockenable2;
  wire             descriptor_memory_s1_unreg_firsttransfer;
  wire             descriptor_memory_s1_waits_for_read;
  wire             descriptor_memory_s1_waits_for_write;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_descriptor_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1;
  wire             p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_rx_descriptor_read_arbiterlock;
  wire             sgdma_rx_descriptor_read_arbiterlock2;
  wire             sgdma_rx_descriptor_read_continuerequest;
  wire             sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  reg              sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_arbiterlock;
  wire             sgdma_rx_descriptor_write_arbiterlock2;
  wire             sgdma_rx_descriptor_write_continuerequest;
  wire             sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_arbiterlock;
  wire             sgdma_tx_descriptor_read_arbiterlock2;
  wire             sgdma_tx_descriptor_read_continuerequest;
  wire             sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  reg              sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_arbiterlock;
  wire             sgdma_tx_descriptor_write_arbiterlock2;
  wire             sgdma_tx_descriptor_write_continuerequest;
  wire             sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1;
  wire    [ 30: 0] shifted_address_to_descriptor_memory_s1_from_cpu_data_master;
  wire    [ 30: 0] shifted_address_to_descriptor_memory_s1_from_cpu_instruction_master;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write;
  wire             wait_for_descriptor_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~descriptor_memory_s1_end_xfer;
    end


  assign descriptor_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_descriptor_memory_s1 | cpu_instruction_master_qualified_request_descriptor_memory_s1 | sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1));
  //assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata;

  assign cpu_data_master_requests_descriptor_memory_s1 = ({cpu_data_master_address_to_slave[30 : 11] , 11'b0} == 31'h48111800) & (cpu_data_master_read | cpu_data_master_write);
  //descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  assign descriptor_memory_s1_arb_share_set_values = 1;

  //descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign descriptor_memory_s1_non_bursting_master_requests = cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    cpu_instruction_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1;

  //descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign descriptor_memory_s1_any_bursting_master_saved_grant = 0;

  //descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign descriptor_memory_s1_arb_share_counter_next_value = descriptor_memory_s1_firsttransfer ? (descriptor_memory_s1_arb_share_set_values - 1) : |descriptor_memory_s1_arb_share_counter ? (descriptor_memory_s1_arb_share_counter - 1) : 0;

  //descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  assign descriptor_memory_s1_allgrants = (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector);

  //descriptor_memory_s1_end_xfer assignment, which is an e_assign
  assign descriptor_memory_s1_end_xfer = ~(descriptor_memory_s1_waits_for_read | descriptor_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_descriptor_memory_s1 = descriptor_memory_s1_end_xfer & (~descriptor_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign descriptor_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_descriptor_memory_s1 & descriptor_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests);

  //descriptor_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_share_counter <= 0;
      else if (descriptor_memory_s1_arb_counter_enable)
          descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
    end


  //descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_slavearbiterlockenable <= 0;
      else if ((|descriptor_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_descriptor_memory_s1) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests))
          descriptor_memory_s1_slavearbiterlockenable <= |descriptor_memory_s1_arb_share_counter_next_value;
    end


  //cpu/data_master descriptor_memory/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign descriptor_memory_s1_slavearbiterlockenable2 = |descriptor_memory_s1_arb_share_counter_next_value;

  //cpu/data_master descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master descriptor_memory/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 <= cpu_instruction_master_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_descriptor_memory_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = (last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 & cpu_instruction_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 & cpu_instruction_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 & cpu_instruction_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 & cpu_instruction_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_descriptor_memory_s1 & cpu_instruction_master_requests_descriptor_memory_s1);

  //descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign descriptor_memory_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_read_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_read_continuerequest = (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1);

  //sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_write_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_write_continuerequest = (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1);

  //sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_read_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_read_continuerequest = (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1);

  //sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_write_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_write_continuerequest = (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1);

  assign cpu_data_master_qualified_request_descriptor_memory_s1 = cpu_data_master_requests_descriptor_memory_s1 & ~((cpu_data_master_read & ((1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))) | cpu_instruction_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in = cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register = {cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register, cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in};

  //cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid cpu_data_master_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_descriptor_memory_s1 = cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;

  //descriptor_memory_s1_writedata mux, which is an e_mux
  assign descriptor_memory_s1_writedata = (cpu_data_master_granted_descriptor_memory_s1)? cpu_data_master_writedata :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? sgdma_rx_descriptor_write_writedata :
    sgdma_tx_descriptor_write_writedata;

  //mux descriptor_memory_s1_clken, which is an e_mux
  assign descriptor_memory_s1_clken = 1'b1;

  assign cpu_instruction_master_requests_descriptor_memory_s1 = (({cpu_instruction_master_address_to_slave[30 : 11] , 11'b0} == 31'h48111800) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= cpu_data_master_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_descriptor_memory_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1);

  assign cpu_instruction_master_qualified_request_descriptor_memory_s1 = cpu_instruction_master_requests_descriptor_memory_s1 & ~((cpu_instruction_master_read & ((1 < cpu_instruction_master_latency_counter))) | cpu_data_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register_in = cpu_instruction_master_granted_descriptor_memory_s1 & cpu_instruction_master_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register = {cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register, cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register_in};

  //cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register <= p1_cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid cpu_instruction_master_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_descriptor_memory_s1 = cpu_instruction_master_read_data_valid_descriptor_memory_s1_shift_register;

  assign sgdma_rx_descriptor_read_requests_descriptor_memory_s1 = (({sgdma_rx_descriptor_read_address_to_slave[31 : 11] , 11'b0} == 32'h48111800) & (sgdma_rx_descriptor_read_read)) & sgdma_rx_descriptor_read_read;
  assign sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 = sgdma_rx_descriptor_read_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in = sgdma_rx_descriptor_read_granted_descriptor_memory_s1 & sgdma_rx_descriptor_read_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register = {sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register, sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in};

  //sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 = sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;

  assign sgdma_rx_descriptor_write_requests_descriptor_memory_s1 = (({sgdma_rx_descriptor_write_address_to_slave[31 : 11] , 11'b0} == 32'h48111800) & (sgdma_rx_descriptor_write_write)) & sgdma_rx_descriptor_write_write;
  assign sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 = sgdma_rx_descriptor_write_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  assign sgdma_tx_descriptor_read_requests_descriptor_memory_s1 = (({sgdma_tx_descriptor_read_address_to_slave[31 : 11] , 11'b0} == 32'h48111800) & (sgdma_tx_descriptor_read_read)) & sgdma_tx_descriptor_read_read;
  assign sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 = sgdma_tx_descriptor_read_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in = sgdma_tx_descriptor_read_granted_descriptor_memory_s1 & sgdma_tx_descriptor_read_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register = {sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register, sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in};

  //sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 = sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;

  assign sgdma_tx_descriptor_write_requests_descriptor_memory_s1 = (({sgdma_tx_descriptor_write_address_to_slave[31 : 11] , 11'b0} == 32'h48111800) & (sgdma_tx_descriptor_write_write)) & sgdma_tx_descriptor_write_write;
  assign sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 = sgdma_tx_descriptor_write_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock);
  //allow new arb cycle for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock & ~sgdma_rx_descriptor_read_arbiterlock & ~sgdma_rx_descriptor_write_arbiterlock & ~sgdma_tx_descriptor_read_arbiterlock & ~sgdma_tx_descriptor_write_arbiterlock;

  //sgdma_tx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[0] = sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;

  //sgdma_tx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[0];

  //sgdma_tx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[0] && sgdma_tx_descriptor_write_requests_descriptor_memory_s1;

  //sgdma_tx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[1] = sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;

  //sgdma_tx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[1];

  //sgdma_tx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[1] && sgdma_tx_descriptor_read_requests_descriptor_memory_s1;

  //sgdma_rx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[2] = sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;

  //sgdma_rx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[2];

  //sgdma_rx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[2] && sgdma_rx_descriptor_write_requests_descriptor_memory_s1;

  //sgdma_rx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[3] = sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;

  //sgdma_rx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[3];

  //sgdma_rx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[3] && sgdma_rx_descriptor_read_requests_descriptor_memory_s1;

  //cpu/instruction_master assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[4] = cpu_instruction_master_qualified_request_descriptor_memory_s1;

  //cpu/instruction_master grant descriptor_memory/s1, which is an e_assign
  assign cpu_instruction_master_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[4];

  //cpu/instruction_master saved-grant descriptor_memory/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[4] && cpu_instruction_master_requests_descriptor_memory_s1;

  //cpu/data_master assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[5] = cpu_data_master_qualified_request_descriptor_memory_s1;

  //cpu/data_master grant descriptor_memory/s1, which is an e_assign
  assign cpu_data_master_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[5];

  //cpu/data_master saved-grant descriptor_memory/s1, which is an e_assign
  assign cpu_data_master_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[5] && cpu_data_master_requests_descriptor_memory_s1;

  //descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  assign descriptor_memory_s1_chosen_master_double_vector = {descriptor_memory_s1_master_qreq_vector, descriptor_memory_s1_master_qreq_vector} & ({~descriptor_memory_s1_master_qreq_vector, ~descriptor_memory_s1_master_qreq_vector} + descriptor_memory_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign descriptor_memory_s1_arb_winner = (descriptor_memory_s1_allow_new_arb_cycle & | descriptor_memory_s1_grant_vector) ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;

  //saved descriptor_memory_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_saved_chosen_master_vector <= 0;
      else if (descriptor_memory_s1_allow_new_arb_cycle)
          descriptor_memory_s1_saved_chosen_master_vector <= |descriptor_memory_s1_grant_vector ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign descriptor_memory_s1_grant_vector = {(descriptor_memory_s1_chosen_master_double_vector[5] | descriptor_memory_s1_chosen_master_double_vector[11]),
    (descriptor_memory_s1_chosen_master_double_vector[4] | descriptor_memory_s1_chosen_master_double_vector[10]),
    (descriptor_memory_s1_chosen_master_double_vector[3] | descriptor_memory_s1_chosen_master_double_vector[9]),
    (descriptor_memory_s1_chosen_master_double_vector[2] | descriptor_memory_s1_chosen_master_double_vector[8]),
    (descriptor_memory_s1_chosen_master_double_vector[1] | descriptor_memory_s1_chosen_master_double_vector[7]),
    (descriptor_memory_s1_chosen_master_double_vector[0] | descriptor_memory_s1_chosen_master_double_vector[6])};

  //descriptor_memory/s1 chosen master rotated left, which is an e_assign
  assign descriptor_memory_s1_chosen_master_rot_left = (descriptor_memory_s1_arb_winner << 1) ? (descriptor_memory_s1_arb_winner << 1) : 1;

  //descriptor_memory/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_addend <= 1;
      else if (|descriptor_memory_s1_grant_vector)
          descriptor_memory_s1_arb_addend <= descriptor_memory_s1_end_xfer? descriptor_memory_s1_chosen_master_rot_left : descriptor_memory_s1_grant_vector;
    end


  assign descriptor_memory_s1_chipselect = cpu_data_master_granted_descriptor_memory_s1 | cpu_instruction_master_granted_descriptor_memory_s1 | sgdma_rx_descriptor_read_granted_descriptor_memory_s1 | sgdma_rx_descriptor_write_granted_descriptor_memory_s1 | sgdma_tx_descriptor_read_granted_descriptor_memory_s1 | sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  //descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_firsttransfer = descriptor_memory_s1_begins_xfer ? descriptor_memory_s1_unreg_firsttransfer : descriptor_memory_s1_reg_firsttransfer;

  //descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_unreg_firsttransfer = ~(descriptor_memory_s1_slavearbiterlockenable & descriptor_memory_s1_any_continuerequest);

  //descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_reg_firsttransfer <= 1'b1;
      else if (descriptor_memory_s1_begins_xfer)
          descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
    end


  //descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign descriptor_memory_s1_beginbursttransfer_internal = descriptor_memory_s1_begins_xfer;

  //descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign descriptor_memory_s1_arbitration_holdoff_internal = descriptor_memory_s1_begins_xfer & descriptor_memory_s1_firsttransfer;

  //descriptor_memory_s1_write assignment, which is an e_mux
  assign descriptor_memory_s1_write = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_write) | (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  assign shifted_address_to_descriptor_memory_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //descriptor_memory_s1_address mux, which is an e_mux
  assign descriptor_memory_s1_address = (cpu_data_master_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_cpu_data_master >> 2) :
    (cpu_instruction_master_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_cpu_instruction_master >> 2) :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read >> 2) :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write >> 2) :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read >> 2) :
    (shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write >> 2);

  assign shifted_address_to_descriptor_memory_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read = sgdma_rx_descriptor_read_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write = sgdma_rx_descriptor_write_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read = sgdma_tx_descriptor_read_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write = sgdma_tx_descriptor_write_address_to_slave;
  //d1_descriptor_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_descriptor_memory_s1_end_xfer <= 1;
      else 
        d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end


  //descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_read = descriptor_memory_s1_in_a_read_cycle & 0;

  //descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_read_cycle = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_descriptor_memory_s1 & cpu_instruction_master_read) | (sgdma_rx_descriptor_read_granted_descriptor_memory_s1 & sgdma_rx_descriptor_read_read) | (sgdma_tx_descriptor_read_granted_descriptor_memory_s1 & sgdma_tx_descriptor_read_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = descriptor_memory_s1_in_a_read_cycle;

  //descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_write = descriptor_memory_s1_in_a_write_cycle & 0;

  //descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_write_cycle = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_write) | (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = descriptor_memory_s1_in_a_write_cycle;

  assign wait_for_descriptor_memory_s1_counter = 0;
  //descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign descriptor_memory_s1_byteenable = (cpu_data_master_granted_descriptor_memory_s1)? cpu_data_master_byteenable :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? {4 {1'b1}} :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? {4 {1'b1}} :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //descriptor_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_descriptor_memory_s1 + cpu_instruction_master_granted_descriptor_memory_s1 + sgdma_rx_descriptor_read_granted_descriptor_memory_s1 + sgdma_rx_descriptor_write_granted_descriptor_memory_s1 + sgdma_tx_descriptor_read_granted_descriptor_memory_s1 + sgdma_tx_descriptor_write_granted_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_descriptor_memory_s1 + cpu_instruction_master_saved_grant_descriptor_memory_s1 + sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 + sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 + sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 + sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_tristate_bridge_avalon_slave_arbitrator (
                                                       // inputs:
                                                        clk,
                                                        cpu_data_master_address_to_slave,
                                                        cpu_data_master_byteenable,
                                                        cpu_data_master_dbs_address,
                                                        cpu_data_master_dbs_write_16,
                                                        cpu_data_master_latency_counter,
                                                        cpu_data_master_read,
                                                        cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                                        cpu_data_master_write,
                                                        cpu_instruction_master_address_to_slave,
                                                        cpu_instruction_master_dbs_address,
                                                        cpu_instruction_master_latency_counter,
                                                        cpu_instruction_master_read,
                                                        reset_n,

                                                       // outputs:
                                                        cpu_data_master_byteenable_ext_flash_s1,
                                                        cpu_data_master_granted_ext_flash_s1,
                                                        cpu_data_master_qualified_request_ext_flash_s1,
                                                        cpu_data_master_read_data_valid_ext_flash_s1,
                                                        cpu_data_master_requests_ext_flash_s1,
                                                        cpu_instruction_master_granted_ext_flash_s1,
                                                        cpu_instruction_master_qualified_request_ext_flash_s1,
                                                        cpu_instruction_master_read_data_valid_ext_flash_s1,
                                                        cpu_instruction_master_requests_ext_flash_s1,
                                                        d1_flash_tristate_bridge_avalon_slave_end_xfer,
                                                        ext_flash_s1_wait_counter_eq_0,
                                                        flash_tristate_bridge_address,
                                                        flash_tristate_bridge_data,
                                                        flash_tristate_bridge_readn,
                                                        flash_tristate_bridge_writen,
                                                        incoming_flash_tristate_bridge_data,
                                                        incoming_flash_tristate_bridge_data_with_Xs_converted_to_0,
                                                        select_n_to_the_ext_flash
                                                     )
;

  output  [  1: 0] cpu_data_master_byteenable_ext_flash_s1;
  output           cpu_data_master_granted_ext_flash_s1;
  output           cpu_data_master_qualified_request_ext_flash_s1;
  output           cpu_data_master_read_data_valid_ext_flash_s1;
  output           cpu_data_master_requests_ext_flash_s1;
  output           cpu_instruction_master_granted_ext_flash_s1;
  output           cpu_instruction_master_qualified_request_ext_flash_s1;
  output           cpu_instruction_master_read_data_valid_ext_flash_s1;
  output           cpu_instruction_master_requests_ext_flash_s1;
  output           d1_flash_tristate_bridge_avalon_slave_end_xfer;
  output           ext_flash_s1_wait_counter_eq_0;
  output  [ 25: 0] flash_tristate_bridge_address;
  inout   [ 15: 0] flash_tristate_bridge_data;
  output           flash_tristate_bridge_readn;
  output           flash_tristate_bridge_writen;
  output  [ 15: 0] incoming_flash_tristate_bridge_data;
  output  [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  output           select_n_to_the_ext_flash;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_dbs_address;
  input   [ 15: 0] cpu_data_master_dbs_write_16;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 30: 0] cpu_instruction_master_address_to_slave;
  input   [  1: 0] cpu_instruction_master_dbs_address;
  input   [  1: 0] cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire    [  1: 0] cpu_data_master_byteenable_ext_flash_s1;
  wire    [  1: 0] cpu_data_master_byteenable_ext_flash_s1_segment_0;
  wire    [  1: 0] cpu_data_master_byteenable_ext_flash_s1_segment_1;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_ext_flash_s1;
  wire             cpu_data_master_qualified_request_ext_flash_s1;
  wire             cpu_data_master_read_data_valid_ext_flash_s1;
  reg     [  1: 0] cpu_data_master_read_data_valid_ext_flash_s1_shift_register;
  wire             cpu_data_master_read_data_valid_ext_flash_s1_shift_register_in;
  wire             cpu_data_master_requests_ext_flash_s1;
  wire             cpu_data_master_saved_grant_ext_flash_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_ext_flash_s1;
  wire             cpu_instruction_master_qualified_request_ext_flash_s1;
  wire             cpu_instruction_master_read_data_valid_ext_flash_s1;
  reg     [  1: 0] cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register;
  wire             cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register_in;
  wire             cpu_instruction_master_requests_ext_flash_s1;
  wire             cpu_instruction_master_saved_grant_ext_flash_s1;
  reg              d1_flash_tristate_bridge_avalon_slave_end_xfer;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 15: 0] d1_outgoing_flash_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave;
  wire    [  5: 0] ext_flash_s1_counter_load_value;
  wire             ext_flash_s1_in_a_read_cycle;
  wire             ext_flash_s1_in_a_write_cycle;
  reg     [  5: 0] ext_flash_s1_wait_counter;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire             ext_flash_s1_waits_for_read;
  wire             ext_flash_s1_waits_for_write;
  wire             ext_flash_s1_with_write_latency;
  reg     [ 25: 0] flash_tristate_bridge_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             flash_tristate_bridge_avalon_slave_allgrants;
  wire             flash_tristate_bridge_avalon_slave_allow_new_arb_cycle;
  wire             flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant;
  wire             flash_tristate_bridge_avalon_slave_any_continuerequest;
  reg     [  1: 0] flash_tristate_bridge_avalon_slave_arb_addend;
  wire             flash_tristate_bridge_avalon_slave_arb_counter_enable;
  reg     [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_counter;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_set_values;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_arb_winner;
  wire             flash_tristate_bridge_avalon_slave_arbitration_holdoff_internal;
  wire             flash_tristate_bridge_avalon_slave_beginbursttransfer_internal;
  wire             flash_tristate_bridge_avalon_slave_begins_xfer;
  wire    [  3: 0] flash_tristate_bridge_avalon_slave_chosen_master_double_vector;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_chosen_master_rot_left;
  wire             flash_tristate_bridge_avalon_slave_end_xfer;
  wire             flash_tristate_bridge_avalon_slave_firsttransfer;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_grant_vector;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_master_qreq_vector;
  wire             flash_tristate_bridge_avalon_slave_non_bursting_master_requests;
  wire             flash_tristate_bridge_avalon_slave_read_pending;
  reg              flash_tristate_bridge_avalon_slave_reg_firsttransfer;
  reg     [  1: 0] flash_tristate_bridge_avalon_slave_saved_chosen_master_vector;
  reg              flash_tristate_bridge_avalon_slave_slavearbiterlockenable;
  wire             flash_tristate_bridge_avalon_slave_slavearbiterlockenable2;
  wire             flash_tristate_bridge_avalon_slave_unreg_firsttransfer;
  wire             flash_tristate_bridge_avalon_slave_write_pending;
  wire    [ 15: 0] flash_tristate_bridge_data;
  reg              flash_tristate_bridge_readn /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              flash_tristate_bridge_writen /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 15: 0] incoming_flash_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_flash_tristate_bridge_data_bit_0_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_10_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_11_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_12_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_13_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_14_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_15_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_1_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_2_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_3_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_4_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_5_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_6_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_7_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_8_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_9_is_x;
  wire    [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  reg              last_cycle_cpu_data_master_granted_slave_ext_flash_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_ext_flash_s1;
  wire    [ 15: 0] outgoing_flash_tristate_bridge_data;
  wire    [  1: 0] p1_cpu_data_master_read_data_valid_ext_flash_s1_shift_register;
  wire    [  1: 0] p1_cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register;
  wire    [ 25: 0] p1_flash_tristate_bridge_address;
  wire             p1_flash_tristate_bridge_readn;
  wire             p1_flash_tristate_bridge_writen;
  wire             p1_select_n_to_the_ext_flash;
  reg              select_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             time_to_write;
  wire             wait_for_ext_flash_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~flash_tristate_bridge_avalon_slave_end_xfer;
    end


  assign flash_tristate_bridge_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_ext_flash_s1 | cpu_instruction_master_qualified_request_ext_flash_s1));
  assign cpu_data_master_requests_ext_flash_s1 = ({cpu_data_master_address_to_slave[30 : 26] , 26'b0} == 31'h44000000) & (cpu_data_master_read | cpu_data_master_write);
  //~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_flash <= ~0;
      else 
        select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end


  assign flash_tristate_bridge_avalon_slave_write_pending = 0;
  //flash_tristate_bridge/avalon_slave read pending calc, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_read_pending = 0;

  //flash_tristate_bridge_avalon_slave_arb_share_counter set values, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_arb_share_set_values = (cpu_data_master_granted_ext_flash_s1)? 2 :
    (cpu_instruction_master_granted_ext_flash_s1)? 2 :
    (cpu_data_master_granted_ext_flash_s1)? 2 :
    (cpu_instruction_master_granted_ext_flash_s1)? 2 :
    1;

  //flash_tristate_bridge_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_non_bursting_master_requests = cpu_data_master_requests_ext_flash_s1 |
    cpu_instruction_master_requests_ext_flash_s1 |
    cpu_data_master_requests_ext_flash_s1 |
    cpu_instruction_master_requests_ext_flash_s1;

  //flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant = 0;

  //flash_tristate_bridge_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_arb_share_counter_next_value = flash_tristate_bridge_avalon_slave_firsttransfer ? (flash_tristate_bridge_avalon_slave_arb_share_set_values - 1) : |flash_tristate_bridge_avalon_slave_arb_share_counter ? (flash_tristate_bridge_avalon_slave_arb_share_counter - 1) : 0;

  //flash_tristate_bridge_avalon_slave_allgrants all slave grants, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_allgrants = (|flash_tristate_bridge_avalon_slave_grant_vector) |
    (|flash_tristate_bridge_avalon_slave_grant_vector) |
    (|flash_tristate_bridge_avalon_slave_grant_vector) |
    (|flash_tristate_bridge_avalon_slave_grant_vector);

  //flash_tristate_bridge_avalon_slave_end_xfer assignment, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_end_xfer = ~(ext_flash_s1_waits_for_read | ext_flash_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave = flash_tristate_bridge_avalon_slave_end_xfer & (~flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //flash_tristate_bridge_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & flash_tristate_bridge_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & ~flash_tristate_bridge_avalon_slave_non_bursting_master_requests);

  //flash_tristate_bridge_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_arb_share_counter <= 0;
      else if (flash_tristate_bridge_avalon_slave_arb_counter_enable)
          flash_tristate_bridge_avalon_slave_arb_share_counter <= flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //flash_tristate_bridge_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|flash_tristate_bridge_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave) | (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & ~flash_tristate_bridge_avalon_slave_non_bursting_master_requests))
          flash_tristate_bridge_avalon_slave_slavearbiterlockenable <= |flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //cpu/data_master flash_tristate_bridge/avalon_slave arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = flash_tristate_bridge_avalon_slave_slavearbiterlockenable & cpu_data_master_continuerequest;

  //flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 = |flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;

  //cpu/data_master flash_tristate_bridge/avalon_slave arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master flash_tristate_bridge/avalon_slave arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = flash_tristate_bridge_avalon_slave_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master flash_tristate_bridge/avalon_slave arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted ext_flash/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_ext_flash_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_ext_flash_s1 <= cpu_instruction_master_saved_grant_ext_flash_s1 ? 1 : (flash_tristate_bridge_avalon_slave_arbitration_holdoff_internal | ~cpu_instruction_master_requests_ext_flash_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_ext_flash_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_ext_flash_s1 & cpu_instruction_master_requests_ext_flash_s1;

  //flash_tristate_bridge_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_ext_flash_s1 = cpu_data_master_requests_ext_flash_s1 & ~((cpu_data_master_read & (flash_tristate_bridge_avalon_slave_write_pending | (flash_tristate_bridge_avalon_slave_read_pending) | (2 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))) | ((flash_tristate_bridge_avalon_slave_read_pending | !cpu_data_master_byteenable_ext_flash_s1) & cpu_data_master_write) | cpu_instruction_master_arbiterlock);
  //cpu_data_master_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_data_master_read_data_valid_ext_flash_s1_shift_register_in = cpu_data_master_granted_ext_flash_s1 & cpu_data_master_read & ~ext_flash_s1_waits_for_read;

  //shift register p1 cpu_data_master_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_data_master_read_data_valid_ext_flash_s1_shift_register = {cpu_data_master_read_data_valid_ext_flash_s1_shift_register, cpu_data_master_read_data_valid_ext_flash_s1_shift_register_in};

  //cpu_data_master_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_data_valid_ext_flash_s1_shift_register <= 0;
      else 
        cpu_data_master_read_data_valid_ext_flash_s1_shift_register <= p1_cpu_data_master_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid cpu_data_master_read_data_valid_ext_flash_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_ext_flash_s1 = cpu_data_master_read_data_valid_ext_flash_s1_shift_register[1];

  //flash_tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_flash_tristate_bridge_data <= 0;
      else 
        incoming_flash_tristate_bridge_data <= flash_tristate_bridge_data;
    end


  //ext_flash_s1_with_write_latency assignment, which is an e_assign
  assign ext_flash_s1_with_write_latency = in_a_write_cycle & (cpu_data_master_qualified_request_ext_flash_s1 | cpu_instruction_master_qualified_request_ext_flash_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (ext_flash_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_flash_tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_flash_tristate_bridge_data <= 0;
      else 
        d1_outgoing_flash_tristate_bridge_data <= outgoing_flash_tristate_bridge_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_flash_tristate_bridge_data tristate driver, which is an e_assign
  assign flash_tristate_bridge_data = (d1_in_a_write_cycle)? d1_outgoing_flash_tristate_bridge_data:{16{1'bz}};

  //outgoing_flash_tristate_bridge_data mux, which is an e_mux
  assign outgoing_flash_tristate_bridge_data = cpu_data_master_dbs_write_16;

  assign cpu_instruction_master_requests_ext_flash_s1 = (({cpu_instruction_master_address_to_slave[30 : 26] , 26'b0} == 31'h44000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted ext_flash/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_ext_flash_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_ext_flash_s1 <= cpu_data_master_saved_grant_ext_flash_s1 ? 1 : (flash_tristate_bridge_avalon_slave_arbitration_holdoff_internal | ~cpu_data_master_requests_ext_flash_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_ext_flash_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_ext_flash_s1 & cpu_data_master_requests_ext_flash_s1;

  assign cpu_instruction_master_qualified_request_ext_flash_s1 = cpu_instruction_master_requests_ext_flash_s1 & ~((cpu_instruction_master_read & (flash_tristate_bridge_avalon_slave_write_pending | (flash_tristate_bridge_avalon_slave_read_pending) | (2 < cpu_instruction_master_latency_counter))) | cpu_data_master_arbiterlock);
  //cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register_in = cpu_instruction_master_granted_ext_flash_s1 & cpu_instruction_master_read & ~ext_flash_s1_waits_for_read;

  //shift register p1 cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register = {cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register, cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register_in};

  //cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register <= 0;
      else 
        cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register <= p1_cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid cpu_instruction_master_read_data_valid_ext_flash_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_ext_flash_s1 = cpu_instruction_master_read_data_valid_ext_flash_s1_shift_register[1];

  //allow new arb cycle for flash_tristate_bridge/avalon_slave, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_master_qreq_vector[0] = cpu_instruction_master_qualified_request_ext_flash_s1;

  //cpu/instruction_master grant ext_flash/s1, which is an e_assign
  assign cpu_instruction_master_granted_ext_flash_s1 = flash_tristate_bridge_avalon_slave_grant_vector[0];

  //cpu/instruction_master saved-grant ext_flash/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_ext_flash_s1 = flash_tristate_bridge_avalon_slave_arb_winner[0] && cpu_instruction_master_requests_ext_flash_s1;

  //cpu/data_master assignment into master qualified-requests vector for ext_flash/s1, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_master_qreq_vector[1] = cpu_data_master_qualified_request_ext_flash_s1;

  //cpu/data_master grant ext_flash/s1, which is an e_assign
  assign cpu_data_master_granted_ext_flash_s1 = flash_tristate_bridge_avalon_slave_grant_vector[1];

  //cpu/data_master saved-grant ext_flash/s1, which is an e_assign
  assign cpu_data_master_saved_grant_ext_flash_s1 = flash_tristate_bridge_avalon_slave_arb_winner[1] && cpu_data_master_requests_ext_flash_s1;

  //flash_tristate_bridge/avalon_slave chosen-master double-vector, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_chosen_master_double_vector = {flash_tristate_bridge_avalon_slave_master_qreq_vector, flash_tristate_bridge_avalon_slave_master_qreq_vector} & ({~flash_tristate_bridge_avalon_slave_master_qreq_vector, ~flash_tristate_bridge_avalon_slave_master_qreq_vector} + flash_tristate_bridge_avalon_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign flash_tristate_bridge_avalon_slave_arb_winner = (flash_tristate_bridge_avalon_slave_allow_new_arb_cycle & | flash_tristate_bridge_avalon_slave_grant_vector) ? flash_tristate_bridge_avalon_slave_grant_vector : flash_tristate_bridge_avalon_slave_saved_chosen_master_vector;

  //saved flash_tristate_bridge_avalon_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_saved_chosen_master_vector <= 0;
      else if (flash_tristate_bridge_avalon_slave_allow_new_arb_cycle)
          flash_tristate_bridge_avalon_slave_saved_chosen_master_vector <= |flash_tristate_bridge_avalon_slave_grant_vector ? flash_tristate_bridge_avalon_slave_grant_vector : flash_tristate_bridge_avalon_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign flash_tristate_bridge_avalon_slave_grant_vector = {(flash_tristate_bridge_avalon_slave_chosen_master_double_vector[1] | flash_tristate_bridge_avalon_slave_chosen_master_double_vector[3]),
    (flash_tristate_bridge_avalon_slave_chosen_master_double_vector[0] | flash_tristate_bridge_avalon_slave_chosen_master_double_vector[2])};

  //flash_tristate_bridge/avalon_slave chosen master rotated left, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_chosen_master_rot_left = (flash_tristate_bridge_avalon_slave_arb_winner << 1) ? (flash_tristate_bridge_avalon_slave_arb_winner << 1) : 1;

  //flash_tristate_bridge/avalon_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_arb_addend <= 1;
      else if (|flash_tristate_bridge_avalon_slave_grant_vector)
          flash_tristate_bridge_avalon_slave_arb_addend <= flash_tristate_bridge_avalon_slave_end_xfer? flash_tristate_bridge_avalon_slave_chosen_master_rot_left : flash_tristate_bridge_avalon_slave_grant_vector;
    end


  assign p1_select_n_to_the_ext_flash = ~(cpu_data_master_granted_ext_flash_s1 | cpu_instruction_master_granted_ext_flash_s1);
  //flash_tristate_bridge_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_firsttransfer = flash_tristate_bridge_avalon_slave_begins_xfer ? flash_tristate_bridge_avalon_slave_unreg_firsttransfer : flash_tristate_bridge_avalon_slave_reg_firsttransfer;

  //flash_tristate_bridge_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_unreg_firsttransfer = ~(flash_tristate_bridge_avalon_slave_slavearbiterlockenable & flash_tristate_bridge_avalon_slave_any_continuerequest);

  //flash_tristate_bridge_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (flash_tristate_bridge_avalon_slave_begins_xfer)
          flash_tristate_bridge_avalon_slave_reg_firsttransfer <= flash_tristate_bridge_avalon_slave_unreg_firsttransfer;
    end


  //flash_tristate_bridge_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_beginbursttransfer_internal = flash_tristate_bridge_avalon_slave_begins_xfer;

  //flash_tristate_bridge_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_arbitration_holdoff_internal = flash_tristate_bridge_avalon_slave_begins_xfer & flash_tristate_bridge_avalon_slave_firsttransfer;

  //~flash_tristate_bridge_readn of type read to ~p1_flash_tristate_bridge_readn, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_readn <= ~0;
      else 
        flash_tristate_bridge_readn <= p1_flash_tristate_bridge_readn;
    end


  //~p1_flash_tristate_bridge_readn assignment, which is an e_mux
  assign p1_flash_tristate_bridge_readn = ~(((cpu_data_master_granted_ext_flash_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_ext_flash_s1 & cpu_instruction_master_read))& ~flash_tristate_bridge_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter < 32));

  //~flash_tristate_bridge_writen of type write to ~p1_flash_tristate_bridge_writen, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_writen <= ~0;
      else 
        flash_tristate_bridge_writen <= p1_flash_tristate_bridge_writen;
    end


  //~p1_flash_tristate_bridge_writen assignment, which is an e_mux
  assign p1_flash_tristate_bridge_writen = ~(((cpu_data_master_granted_ext_flash_s1 & cpu_data_master_write)) & ~flash_tristate_bridge_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter >= 8) & (ext_flash_s1_wait_counter < 40));

  //flash_tristate_bridge_address of type address to p1_flash_tristate_bridge_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_address <= 0;
      else 
        flash_tristate_bridge_address <= p1_flash_tristate_bridge_address;
    end


  //p1_flash_tristate_bridge_address mux, which is an e_mux
  assign p1_flash_tristate_bridge_address = (cpu_data_master_granted_ext_flash_s1)? ({cpu_data_master_address_to_slave >> 2,
    cpu_data_master_dbs_address[1],
    {1 {1'b0}}}) :
    ({cpu_instruction_master_address_to_slave >> 2,
    cpu_instruction_master_dbs_address[1],
    {1 {1'b0}}});

  //d1_flash_tristate_bridge_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_flash_tristate_bridge_avalon_slave_end_xfer <= 1;
      else 
        d1_flash_tristate_bridge_avalon_slave_end_xfer <= flash_tristate_bridge_avalon_slave_end_xfer;
    end


  //ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_read = ext_flash_s1_in_a_read_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_read_cycle = (cpu_data_master_granted_ext_flash_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_ext_flash_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ext_flash_s1_in_a_read_cycle;

  //ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_write = ext_flash_s1_in_a_write_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_write_cycle = cpu_data_master_granted_ext_flash_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ext_flash_s1_in_a_write_cycle;

  assign ext_flash_s1_wait_counter_eq_0 = ext_flash_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_s1_wait_counter <= 0;
      else 
        ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end


  assign ext_flash_s1_counter_load_value = ((ext_flash_s1_in_a_read_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 52 :
    ((ext_flash_s1_in_a_write_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 60 :
    (~ext_flash_s1_wait_counter_eq_0)? ext_flash_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_flash_s1_counter = flash_tristate_bridge_avalon_slave_begins_xfer | ~ext_flash_s1_wait_counter_eq_0;
  assign {cpu_data_master_byteenable_ext_flash_s1_segment_1,
cpu_data_master_byteenable_ext_flash_s1_segment_0} = cpu_data_master_byteenable;
  assign cpu_data_master_byteenable_ext_flash_s1 = ((cpu_data_master_dbs_address[1] == 0))? cpu_data_master_byteenable_ext_flash_s1_segment_0 :
    cpu_data_master_byteenable_ext_flash_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //incoming_flash_tristate_bridge_data_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_0_is_x = ^(incoming_flash_tristate_bridge_data[0]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[0] = incoming_flash_tristate_bridge_data_bit_0_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[0];

  //incoming_flash_tristate_bridge_data_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_1_is_x = ^(incoming_flash_tristate_bridge_data[1]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[1] = incoming_flash_tristate_bridge_data_bit_1_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[1];

  //incoming_flash_tristate_bridge_data_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_2_is_x = ^(incoming_flash_tristate_bridge_data[2]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[2] = incoming_flash_tristate_bridge_data_bit_2_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[2];

  //incoming_flash_tristate_bridge_data_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_3_is_x = ^(incoming_flash_tristate_bridge_data[3]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[3] = incoming_flash_tristate_bridge_data_bit_3_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[3];

  //incoming_flash_tristate_bridge_data_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_4_is_x = ^(incoming_flash_tristate_bridge_data[4]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[4] = incoming_flash_tristate_bridge_data_bit_4_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[4];

  //incoming_flash_tristate_bridge_data_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_5_is_x = ^(incoming_flash_tristate_bridge_data[5]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[5] = incoming_flash_tristate_bridge_data_bit_5_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[5];

  //incoming_flash_tristate_bridge_data_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_6_is_x = ^(incoming_flash_tristate_bridge_data[6]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[6] = incoming_flash_tristate_bridge_data_bit_6_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[6];

  //incoming_flash_tristate_bridge_data_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_7_is_x = ^(incoming_flash_tristate_bridge_data[7]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[7] = incoming_flash_tristate_bridge_data_bit_7_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[7];

  //incoming_flash_tristate_bridge_data_bit_8_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_8_is_x = ^(incoming_flash_tristate_bridge_data[8]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[8] = incoming_flash_tristate_bridge_data_bit_8_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[8];

  //incoming_flash_tristate_bridge_data_bit_9_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_9_is_x = ^(incoming_flash_tristate_bridge_data[9]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[9] = incoming_flash_tristate_bridge_data_bit_9_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[9];

  //incoming_flash_tristate_bridge_data_bit_10_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_10_is_x = ^(incoming_flash_tristate_bridge_data[10]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[10] = incoming_flash_tristate_bridge_data_bit_10_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[10];

  //incoming_flash_tristate_bridge_data_bit_11_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_11_is_x = ^(incoming_flash_tristate_bridge_data[11]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[11] = incoming_flash_tristate_bridge_data_bit_11_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[11];

  //incoming_flash_tristate_bridge_data_bit_12_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_12_is_x = ^(incoming_flash_tristate_bridge_data[12]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[12] = incoming_flash_tristate_bridge_data_bit_12_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[12];

  //incoming_flash_tristate_bridge_data_bit_13_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_13_is_x = ^(incoming_flash_tristate_bridge_data[13]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[13] = incoming_flash_tristate_bridge_data_bit_13_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[13];

  //incoming_flash_tristate_bridge_data_bit_14_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_14_is_x = ^(incoming_flash_tristate_bridge_data[14]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[14] = incoming_flash_tristate_bridge_data_bit_14_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[14];

  //incoming_flash_tristate_bridge_data_bit_15_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_15_is_x = ^(incoming_flash_tristate_bridge_data[15]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15] = incoming_flash_tristate_bridge_data_bit_15_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[15];

  //ext_flash/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_ext_flash_s1 + cpu_instruction_master_granted_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_ext_flash_s1 + cpu_instruction_master_saved_grant_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0 = incoming_flash_tristate_bridge_data;
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_tristate_bridge_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module high_res_timer_s1_arbitrator (
                                      // inputs:
                                       clk,
                                       cpu_data_master_address_to_slave,
                                       cpu_data_master_latency_counter,
                                       cpu_data_master_read,
                                       cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                       cpu_data_master_write,
                                       cpu_data_master_writedata,
                                       high_res_timer_s1_irq,
                                       high_res_timer_s1_readdata,
                                       reset_n,

                                      // outputs:
                                       cpu_data_master_granted_high_res_timer_s1,
                                       cpu_data_master_qualified_request_high_res_timer_s1,
                                       cpu_data_master_read_data_valid_high_res_timer_s1,
                                       cpu_data_master_requests_high_res_timer_s1,
                                       d1_high_res_timer_s1_end_xfer,
                                       high_res_timer_s1_address,
                                       high_res_timer_s1_chipselect,
                                       high_res_timer_s1_irq_from_sa,
                                       high_res_timer_s1_readdata_from_sa,
                                       high_res_timer_s1_reset_n,
                                       high_res_timer_s1_write_n,
                                       high_res_timer_s1_writedata
                                    )
;

  output           cpu_data_master_granted_high_res_timer_s1;
  output           cpu_data_master_qualified_request_high_res_timer_s1;
  output           cpu_data_master_read_data_valid_high_res_timer_s1;
  output           cpu_data_master_requests_high_res_timer_s1;
  output           d1_high_res_timer_s1_end_xfer;
  output  [  2: 0] high_res_timer_s1_address;
  output           high_res_timer_s1_chipselect;
  output           high_res_timer_s1_irq_from_sa;
  output  [ 15: 0] high_res_timer_s1_readdata_from_sa;
  output           high_res_timer_s1_reset_n;
  output           high_res_timer_s1_write_n;
  output  [ 15: 0] high_res_timer_s1_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            high_res_timer_s1_irq;
  input   [ 15: 0] high_res_timer_s1_readdata;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_high_res_timer_s1;
  wire             cpu_data_master_qualified_request_high_res_timer_s1;
  wire             cpu_data_master_read_data_valid_high_res_timer_s1;
  wire             cpu_data_master_requests_high_res_timer_s1;
  wire             cpu_data_master_saved_grant_high_res_timer_s1;
  reg              d1_high_res_timer_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_high_res_timer_s1;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_allgrants;
  wire             high_res_timer_s1_allow_new_arb_cycle;
  wire             high_res_timer_s1_any_bursting_master_saved_grant;
  wire             high_res_timer_s1_any_continuerequest;
  wire             high_res_timer_s1_arb_counter_enable;
  reg     [  1: 0] high_res_timer_s1_arb_share_counter;
  wire    [  1: 0] high_res_timer_s1_arb_share_counter_next_value;
  wire    [  1: 0] high_res_timer_s1_arb_share_set_values;
  wire             high_res_timer_s1_beginbursttransfer_internal;
  wire             high_res_timer_s1_begins_xfer;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_end_xfer;
  wire             high_res_timer_s1_firsttransfer;
  wire             high_res_timer_s1_grant_vector;
  wire             high_res_timer_s1_in_a_read_cycle;
  wire             high_res_timer_s1_in_a_write_cycle;
  wire             high_res_timer_s1_irq_from_sa;
  wire             high_res_timer_s1_master_qreq_vector;
  wire             high_res_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  reg              high_res_timer_s1_reg_firsttransfer;
  wire             high_res_timer_s1_reset_n;
  reg              high_res_timer_s1_slavearbiterlockenable;
  wire             high_res_timer_s1_slavearbiterlockenable2;
  wire             high_res_timer_s1_unreg_firsttransfer;
  wire             high_res_timer_s1_waits_for_read;
  wire             high_res_timer_s1_waits_for_write;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_high_res_timer_s1_from_cpu_data_master;
  wire             wait_for_high_res_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~high_res_timer_s1_end_xfer;
    end


  assign high_res_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_high_res_timer_s1));
  //assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata;

  assign cpu_data_master_requests_high_res_timer_s1 = ({cpu_data_master_address_to_slave[30 : 5] , 5'b0} == 31'h48112500) & (cpu_data_master_read | cpu_data_master_write);
  //high_res_timer_s1_arb_share_counter set values, which is an e_mux
  assign high_res_timer_s1_arb_share_set_values = 1;

  //high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign high_res_timer_s1_non_bursting_master_requests = cpu_data_master_requests_high_res_timer_s1;

  //high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign high_res_timer_s1_any_bursting_master_saved_grant = 0;

  //high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign high_res_timer_s1_arb_share_counter_next_value = high_res_timer_s1_firsttransfer ? (high_res_timer_s1_arb_share_set_values - 1) : |high_res_timer_s1_arb_share_counter ? (high_res_timer_s1_arb_share_counter - 1) : 0;

  //high_res_timer_s1_allgrants all slave grants, which is an e_mux
  assign high_res_timer_s1_allgrants = |high_res_timer_s1_grant_vector;

  //high_res_timer_s1_end_xfer assignment, which is an e_assign
  assign high_res_timer_s1_end_xfer = ~(high_res_timer_s1_waits_for_read | high_res_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_high_res_timer_s1 = high_res_timer_s1_end_xfer & (~high_res_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign high_res_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_high_res_timer_s1 & high_res_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests);

  //high_res_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_arb_share_counter <= 0;
      else if (high_res_timer_s1_arb_counter_enable)
          high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
    end


  //high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_slavearbiterlockenable <= 0;
      else if ((|high_res_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_high_res_timer_s1) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests))
          high_res_timer_s1_slavearbiterlockenable <= |high_res_timer_s1_arb_share_counter_next_value;
    end


  //cpu/data_master high_res_timer/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = high_res_timer_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign high_res_timer_s1_slavearbiterlockenable2 = |high_res_timer_s1_arb_share_counter_next_value;

  //cpu/data_master high_res_timer/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = high_res_timer_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign high_res_timer_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_high_res_timer_s1 = cpu_data_master_requests_high_res_timer_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_high_res_timer_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_high_res_timer_s1 = cpu_data_master_granted_high_res_timer_s1 & cpu_data_master_read & ~high_res_timer_s1_waits_for_read;

  //high_res_timer_s1_writedata mux, which is an e_mux
  assign high_res_timer_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_high_res_timer_s1 = cpu_data_master_qualified_request_high_res_timer_s1;

  //cpu/data_master saved-grant high_res_timer/s1, which is an e_assign
  assign cpu_data_master_saved_grant_high_res_timer_s1 = cpu_data_master_requests_high_res_timer_s1;

  //allow new arb cycle for high_res_timer/s1, which is an e_assign
  assign high_res_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign high_res_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign high_res_timer_s1_master_qreq_vector = 1;

  //high_res_timer_s1_reset_n assignment, which is an e_assign
  assign high_res_timer_s1_reset_n = reset_n;

  assign high_res_timer_s1_chipselect = cpu_data_master_granted_high_res_timer_s1;
  //high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_firsttransfer = high_res_timer_s1_begins_xfer ? high_res_timer_s1_unreg_firsttransfer : high_res_timer_s1_reg_firsttransfer;

  //high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_unreg_firsttransfer = ~(high_res_timer_s1_slavearbiterlockenable & high_res_timer_s1_any_continuerequest);

  //high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_reg_firsttransfer <= 1'b1;
      else if (high_res_timer_s1_begins_xfer)
          high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
    end


  //high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign high_res_timer_s1_beginbursttransfer_internal = high_res_timer_s1_begins_xfer;

  //~high_res_timer_s1_write_n assignment, which is an e_mux
  assign high_res_timer_s1_write_n = ~(cpu_data_master_granted_high_res_timer_s1 & cpu_data_master_write);

  assign shifted_address_to_high_res_timer_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //high_res_timer_s1_address mux, which is an e_mux
  assign high_res_timer_s1_address = shifted_address_to_high_res_timer_s1_from_cpu_data_master >> 2;

  //d1_high_res_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_high_res_timer_s1_end_xfer <= 1;
      else 
        d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end


  //high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_read = high_res_timer_s1_in_a_read_cycle & high_res_timer_s1_begins_xfer;

  //high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_read_cycle = cpu_data_master_granted_high_res_timer_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = high_res_timer_s1_in_a_read_cycle;

  //high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_write = high_res_timer_s1_in_a_write_cycle & 0;

  //high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_write_cycle = cpu_data_master_granted_high_res_timer_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = high_res_timer_s1_in_a_write_cycle;

  assign wait_for_high_res_timer_s1_counter = 0;
  //assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //high_res_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_data_master_address_to_slave,
                                                 cpu_data_master_latency_counter,
                                                 cpu_data_master_read,
                                                 cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                                 cpu_data_master_write,
                                                 cpu_data_master_writedata,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata
                                              )
;

  output           cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave;
  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg     [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire    [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  1: 0] jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire    [ 30: 0] shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign cpu_data_master_requests_jtag_uart_avalon_jtag_slave = ({cpu_data_master_address_to_slave[30 : 3] , 3'b0} == 31'h48112840) & (cpu_data_master_read | cpu_data_master_write);
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = cpu_data_master_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & cpu_data_master_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave = cpu_data_master_requests_jtag_uart_avalon_jtag_slave & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave = cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_read & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_jtag_uart_avalon_jtag_slave = cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;

  //cpu/data_master saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave = cpu_data_master_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_read);

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_write);

  assign shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master = cpu_data_master_address_to_slave;
  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master >> 2;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = cpu_data_master_granted_jtag_uart_avalon_jtag_slave & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module master_read_avalon_master_arbitrator (
                                              // inputs:
                                               clk,
                                               clock_crossing_master_ddr2_s1_readdata_from_sa,
                                               clock_crossing_master_ddr2_s1_waitrequest_from_sa,
                                               d1_clock_crossing_master_ddr2_s1_end_xfer,
                                               master_read_avalon_master_address,
                                               master_read_avalon_master_burstcount,
                                               master_read_avalon_master_byteenable,
                                               master_read_avalon_master_read,
                                               master_read_granted_clock_crossing_master_ddr2_s1,
                                               master_read_qualified_request_clock_crossing_master_ddr2_s1,
                                               master_read_read_data_valid_clock_crossing_master_ddr2_s1,
                                               master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register,
                                               master_read_requests_clock_crossing_master_ddr2_s1,
                                               reset_n,

                                              // outputs:
                                               master_read_avalon_master_address_to_slave,
                                               master_read_avalon_master_readdata,
                                               master_read_avalon_master_readdatavalid,
                                               master_read_avalon_master_reset,
                                               master_read_avalon_master_waitrequest,
                                               master_read_latency_counter
                                            )
;

  output  [ 29: 0] master_read_avalon_master_address_to_slave;
  output  [255: 0] master_read_avalon_master_readdata;
  output           master_read_avalon_master_readdatavalid;
  output           master_read_avalon_master_reset;
  output           master_read_avalon_master_waitrequest;
  output           master_read_latency_counter;
  input            clk;
  input   [255: 0] clock_crossing_master_ddr2_s1_readdata_from_sa;
  input            clock_crossing_master_ddr2_s1_waitrequest_from_sa;
  input            d1_clock_crossing_master_ddr2_s1_end_xfer;
  input   [ 29: 0] master_read_avalon_master_address;
  input   [  3: 0] master_read_avalon_master_burstcount;
  input   [ 31: 0] master_read_avalon_master_byteenable;
  input            master_read_avalon_master_read;
  input            master_read_granted_clock_crossing_master_ddr2_s1;
  input            master_read_qualified_request_clock_crossing_master_ddr2_s1;
  input            master_read_read_data_valid_clock_crossing_master_ddr2_s1;
  input            master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register;
  input            master_read_requests_clock_crossing_master_ddr2_s1;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  reg     [ 29: 0] master_read_avalon_master_address_last_time;
  wire    [ 29: 0] master_read_avalon_master_address_to_slave;
  reg     [  3: 0] master_read_avalon_master_burstcount_last_time;
  reg     [ 31: 0] master_read_avalon_master_byteenable_last_time;
  wire             master_read_avalon_master_is_granted_some_slave;
  reg              master_read_avalon_master_read_but_no_slave_selected;
  reg              master_read_avalon_master_read_last_time;
  wire    [255: 0] master_read_avalon_master_readdata;
  wire             master_read_avalon_master_readdatavalid;
  wire             master_read_avalon_master_reset;
  wire             master_read_avalon_master_run;
  wire             master_read_avalon_master_waitrequest;
  reg              master_read_latency_counter;
  wire             p1_master_read_latency_counter;
  wire             pre_flush_master_read_avalon_master_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (master_read_qualified_request_clock_crossing_master_ddr2_s1 | ~master_read_requests_clock_crossing_master_ddr2_s1) & (master_read_granted_clock_crossing_master_ddr2_s1 | ~master_read_qualified_request_clock_crossing_master_ddr2_s1) & ((~master_read_qualified_request_clock_crossing_master_ddr2_s1 | ~(master_read_avalon_master_read) | (1 & ~clock_crossing_master_ddr2_s1_waitrequest_from_sa & (master_read_avalon_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign master_read_avalon_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign master_read_avalon_master_address_to_slave = master_read_avalon_master_address[29 : 0];

  //master_read_avalon_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_avalon_master_read_but_no_slave_selected <= 0;
      else 
        master_read_avalon_master_read_but_no_slave_selected <= master_read_avalon_master_read & master_read_avalon_master_run & ~master_read_avalon_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign master_read_avalon_master_is_granted_some_slave = master_read_granted_clock_crossing_master_ddr2_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_master_read_avalon_master_readdatavalid = master_read_read_data_valid_clock_crossing_master_ddr2_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign master_read_avalon_master_readdatavalid = master_read_avalon_master_read_but_no_slave_selected |
    pre_flush_master_read_avalon_master_readdatavalid;

  //master_read/avalon_master readdata mux, which is an e_mux
  assign master_read_avalon_master_readdata = clock_crossing_master_ddr2_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign master_read_avalon_master_waitrequest = ~master_read_avalon_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_latency_counter <= 0;
      else 
        master_read_latency_counter <= p1_master_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_master_read_latency_counter = ((master_read_avalon_master_run & master_read_avalon_master_read))? latency_load_value :
    (master_read_latency_counter)? master_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //~master_read_avalon_master_reset assignment, which is an e_assign
  assign master_read_avalon_master_reset = ~reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //master_read_avalon_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_avalon_master_address_last_time <= 0;
      else 
        master_read_avalon_master_address_last_time <= master_read_avalon_master_address;
    end


  //master_read/avalon_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= master_read_avalon_master_waitrequest & (master_read_avalon_master_read);
    end


  //master_read_avalon_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_read_avalon_master_address != master_read_avalon_master_address_last_time))
        begin
          $write("%0d ns: master_read_avalon_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_read_avalon_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_avalon_master_burstcount_last_time <= 0;
      else 
        master_read_avalon_master_burstcount_last_time <= master_read_avalon_master_burstcount;
    end


  //master_read_avalon_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_read_avalon_master_burstcount != master_read_avalon_master_burstcount_last_time))
        begin
          $write("%0d ns: master_read_avalon_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_read_avalon_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_avalon_master_byteenable_last_time <= 0;
      else 
        master_read_avalon_master_byteenable_last_time <= master_read_avalon_master_byteenable;
    end


  //master_read_avalon_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_read_avalon_master_byteenable != master_read_avalon_master_byteenable_last_time))
        begin
          $write("%0d ns: master_read_avalon_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_read_avalon_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_read_avalon_master_read_last_time <= 0;
      else 
        master_read_avalon_master_read_last_time <= master_read_avalon_master_read;
    end


  //master_read_avalon_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_read_avalon_master_read != master_read_avalon_master_read_last_time))
        begin
          $write("%0d ns: master_read_avalon_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module master_write_avalon_master_arbitrator (
                                               // inputs:
                                                clk,
                                                clock_crossing_master_ddr2_s1_waitrequest_from_sa,
                                                d1_clock_crossing_master_ddr2_s1_end_xfer,
                                                master_write_avalon_master_address,
                                                master_write_avalon_master_burstcount,
                                                master_write_avalon_master_byteenable,
                                                master_write_avalon_master_write,
                                                master_write_avalon_master_writedata,
                                                master_write_granted_clock_crossing_master_ddr2_s1,
                                                master_write_qualified_request_clock_crossing_master_ddr2_s1,
                                                master_write_requests_clock_crossing_master_ddr2_s1,
                                                reset_n,

                                               // outputs:
                                                master_write_avalon_master_address_to_slave,
                                                master_write_avalon_master_reset,
                                                master_write_avalon_master_waitrequest
                                             )
;

  output  [ 29: 0] master_write_avalon_master_address_to_slave;
  output           master_write_avalon_master_reset;
  output           master_write_avalon_master_waitrequest;
  input            clk;
  input            clock_crossing_master_ddr2_s1_waitrequest_from_sa;
  input            d1_clock_crossing_master_ddr2_s1_end_xfer;
  input   [ 29: 0] master_write_avalon_master_address;
  input   [  3: 0] master_write_avalon_master_burstcount;
  input   [ 31: 0] master_write_avalon_master_byteenable;
  input            master_write_avalon_master_write;
  input   [255: 0] master_write_avalon_master_writedata;
  input            master_write_granted_clock_crossing_master_ddr2_s1;
  input            master_write_qualified_request_clock_crossing_master_ddr2_s1;
  input            master_write_requests_clock_crossing_master_ddr2_s1;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 29: 0] master_write_avalon_master_address_last_time;
  wire    [ 29: 0] master_write_avalon_master_address_to_slave;
  reg     [  3: 0] master_write_avalon_master_burstcount_last_time;
  reg     [ 31: 0] master_write_avalon_master_byteenable_last_time;
  wire             master_write_avalon_master_reset;
  wire             master_write_avalon_master_run;
  wire             master_write_avalon_master_waitrequest;
  reg              master_write_avalon_master_write_last_time;
  reg     [255: 0] master_write_avalon_master_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (master_write_qualified_request_clock_crossing_master_ddr2_s1 | ~master_write_requests_clock_crossing_master_ddr2_s1) & (master_write_granted_clock_crossing_master_ddr2_s1 | ~master_write_qualified_request_clock_crossing_master_ddr2_s1) & ((~master_write_qualified_request_clock_crossing_master_ddr2_s1 | ~(master_write_avalon_master_write) | (1 & ~clock_crossing_master_ddr2_s1_waitrequest_from_sa & (master_write_avalon_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign master_write_avalon_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign master_write_avalon_master_address_to_slave = master_write_avalon_master_address[29 : 0];

  //actual waitrequest port, which is an e_assign
  assign master_write_avalon_master_waitrequest = ~master_write_avalon_master_run;

  //~master_write_avalon_master_reset assignment, which is an e_assign
  assign master_write_avalon_master_reset = ~reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //master_write_avalon_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_write_avalon_master_address_last_time <= 0;
      else 
        master_write_avalon_master_address_last_time <= master_write_avalon_master_address;
    end


  //master_write/avalon_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= master_write_avalon_master_waitrequest & (master_write_avalon_master_write);
    end


  //master_write_avalon_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_write_avalon_master_address != master_write_avalon_master_address_last_time))
        begin
          $write("%0d ns: master_write_avalon_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_write_avalon_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_write_avalon_master_burstcount_last_time <= 0;
      else 
        master_write_avalon_master_burstcount_last_time <= master_write_avalon_master_burstcount;
    end


  //master_write_avalon_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_write_avalon_master_burstcount != master_write_avalon_master_burstcount_last_time))
        begin
          $write("%0d ns: master_write_avalon_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_write_avalon_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_write_avalon_master_byteenable_last_time <= 0;
      else 
        master_write_avalon_master_byteenable_last_time <= master_write_avalon_master_byteenable;
    end


  //master_write_avalon_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_write_avalon_master_byteenable != master_write_avalon_master_byteenable_last_time))
        begin
          $write("%0d ns: master_write_avalon_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_write_avalon_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_write_avalon_master_write_last_time <= 0;
      else 
        master_write_avalon_master_write_last_time <= master_write_avalon_master_write;
    end


  //master_write_avalon_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_write_avalon_master_write != master_write_avalon_master_write_last_time))
        begin
          $write("%0d ns: master_write_avalon_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //master_write_avalon_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          master_write_avalon_master_writedata_last_time <= 0;
      else 
        master_write_avalon_master_writedata_last_time <= master_write_avalon_master_writedata;
    end


  //master_write_avalon_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (master_write_avalon_master_writedata != master_write_avalon_master_writedata_last_time) & master_write_avalon_master_write)
        begin
          $write("%0d ns: master_write_avalon_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_memory_s1_arbitrator (
                                     // inputs:
                                      clk,
                                      cpu_data_master_address_to_slave,
                                      cpu_data_master_byteenable,
                                      cpu_data_master_latency_counter,
                                      cpu_data_master_read,
                                      cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                      cpu_data_master_write,
                                      cpu_data_master_writedata,
                                      cpu_instruction_master_address_to_slave,
                                      cpu_instruction_master_latency_counter,
                                      cpu_instruction_master_read,
                                      onchip_memory_s1_readdata,
                                      reset_n,
                                      sgdma_rx_m_write_address_to_slave,
                                      sgdma_rx_m_write_byteenable,
                                      sgdma_rx_m_write_write,
                                      sgdma_rx_m_write_writedata,
                                      sgdma_tx_m_read_address_to_slave,
                                      sgdma_tx_m_read_latency_counter,
                                      sgdma_tx_m_read_read,

                                     // outputs:
                                      cpu_data_master_granted_onchip_memory_s1,
                                      cpu_data_master_qualified_request_onchip_memory_s1,
                                      cpu_data_master_read_data_valid_onchip_memory_s1,
                                      cpu_data_master_requests_onchip_memory_s1,
                                      cpu_instruction_master_granted_onchip_memory_s1,
                                      cpu_instruction_master_qualified_request_onchip_memory_s1,
                                      cpu_instruction_master_read_data_valid_onchip_memory_s1,
                                      cpu_instruction_master_requests_onchip_memory_s1,
                                      d1_onchip_memory_s1_end_xfer,
                                      onchip_memory_s1_address,
                                      onchip_memory_s1_byteenable,
                                      onchip_memory_s1_chipselect,
                                      onchip_memory_s1_clken,
                                      onchip_memory_s1_readdata_from_sa,
                                      onchip_memory_s1_write,
                                      onchip_memory_s1_writedata,
                                      sgdma_rx_m_write_granted_onchip_memory_s1,
                                      sgdma_rx_m_write_qualified_request_onchip_memory_s1,
                                      sgdma_rx_m_write_requests_onchip_memory_s1,
                                      sgdma_tx_m_read_granted_onchip_memory_s1,
                                      sgdma_tx_m_read_qualified_request_onchip_memory_s1,
                                      sgdma_tx_m_read_read_data_valid_onchip_memory_s1,
                                      sgdma_tx_m_read_requests_onchip_memory_s1
                                   )
;

  output           cpu_data_master_granted_onchip_memory_s1;
  output           cpu_data_master_qualified_request_onchip_memory_s1;
  output           cpu_data_master_read_data_valid_onchip_memory_s1;
  output           cpu_data_master_requests_onchip_memory_s1;
  output           cpu_instruction_master_granted_onchip_memory_s1;
  output           cpu_instruction_master_qualified_request_onchip_memory_s1;
  output           cpu_instruction_master_read_data_valid_onchip_memory_s1;
  output           cpu_instruction_master_requests_onchip_memory_s1;
  output           d1_onchip_memory_s1_end_xfer;
  output  [ 16: 0] onchip_memory_s1_address;
  output  [  3: 0] onchip_memory_s1_byteenable;
  output           onchip_memory_s1_chipselect;
  output           onchip_memory_s1_clken;
  output  [ 31: 0] onchip_memory_s1_readdata_from_sa;
  output           onchip_memory_s1_write;
  output  [ 31: 0] onchip_memory_s1_writedata;
  output           sgdma_rx_m_write_granted_onchip_memory_s1;
  output           sgdma_rx_m_write_qualified_request_onchip_memory_s1;
  output           sgdma_rx_m_write_requests_onchip_memory_s1;
  output           sgdma_tx_m_read_granted_onchip_memory_s1;
  output           sgdma_tx_m_read_qualified_request_onchip_memory_s1;
  output           sgdma_tx_m_read_read_data_valid_onchip_memory_s1;
  output           sgdma_tx_m_read_requests_onchip_memory_s1;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 30: 0] cpu_instruction_master_address_to_slave;
  input   [  1: 0] cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input   [ 31: 0] onchip_memory_s1_readdata;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address_to_slave;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;
  input   [ 31: 0] sgdma_tx_m_read_address_to_slave;
  input            sgdma_tx_m_read_latency_counter;
  input            sgdma_tx_m_read_read;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_onchip_memory_s1;
  wire             cpu_data_master_qualified_request_onchip_memory_s1;
  wire             cpu_data_master_read_data_valid_onchip_memory_s1;
  reg              cpu_data_master_read_data_valid_onchip_memory_s1_shift_register;
  wire             cpu_data_master_read_data_valid_onchip_memory_s1_shift_register_in;
  wire             cpu_data_master_requests_onchip_memory_s1;
  wire             cpu_data_master_saved_grant_onchip_memory_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_onchip_memory_s1;
  wire             cpu_instruction_master_qualified_request_onchip_memory_s1;
  wire             cpu_instruction_master_read_data_valid_onchip_memory_s1;
  reg              cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register;
  wire             cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in;
  wire             cpu_instruction_master_requests_onchip_memory_s1;
  wire             cpu_instruction_master_saved_grant_onchip_memory_s1;
  reg              d1_onchip_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_onchip_memory_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1;
  reg              last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1;
  reg              last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1;
  wire    [ 16: 0] onchip_memory_s1_address;
  wire             onchip_memory_s1_allgrants;
  wire             onchip_memory_s1_allow_new_arb_cycle;
  wire             onchip_memory_s1_any_bursting_master_saved_grant;
  wire             onchip_memory_s1_any_continuerequest;
  reg     [  3: 0] onchip_memory_s1_arb_addend;
  wire             onchip_memory_s1_arb_counter_enable;
  reg     [  1: 0] onchip_memory_s1_arb_share_counter;
  wire    [  1: 0] onchip_memory_s1_arb_share_counter_next_value;
  wire    [  1: 0] onchip_memory_s1_arb_share_set_values;
  wire    [  3: 0] onchip_memory_s1_arb_winner;
  wire             onchip_memory_s1_arbitration_holdoff_internal;
  wire             onchip_memory_s1_beginbursttransfer_internal;
  wire             onchip_memory_s1_begins_xfer;
  wire    [  3: 0] onchip_memory_s1_byteenable;
  wire             onchip_memory_s1_chipselect;
  wire    [  7: 0] onchip_memory_s1_chosen_master_double_vector;
  wire    [  3: 0] onchip_memory_s1_chosen_master_rot_left;
  wire             onchip_memory_s1_clken;
  wire             onchip_memory_s1_end_xfer;
  wire             onchip_memory_s1_firsttransfer;
  wire    [  3: 0] onchip_memory_s1_grant_vector;
  wire             onchip_memory_s1_in_a_read_cycle;
  wire             onchip_memory_s1_in_a_write_cycle;
  wire    [  3: 0] onchip_memory_s1_master_qreq_vector;
  wire             onchip_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_memory_s1_readdata_from_sa;
  reg              onchip_memory_s1_reg_firsttransfer;
  reg     [  3: 0] onchip_memory_s1_saved_chosen_master_vector;
  reg              onchip_memory_s1_slavearbiterlockenable;
  wire             onchip_memory_s1_slavearbiterlockenable2;
  wire             onchip_memory_s1_unreg_firsttransfer;
  wire             onchip_memory_s1_waits_for_read;
  wire             onchip_memory_s1_waits_for_write;
  wire             onchip_memory_s1_write;
  wire    [ 31: 0] onchip_memory_s1_writedata;
  wire             p1_cpu_data_master_read_data_valid_onchip_memory_s1_shift_register;
  wire             p1_cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register;
  wire             p1_sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register;
  wire             sgdma_rx_m_write_arbiterlock;
  wire             sgdma_rx_m_write_arbiterlock2;
  wire             sgdma_rx_m_write_continuerequest;
  wire             sgdma_rx_m_write_granted_onchip_memory_s1;
  wire             sgdma_rx_m_write_qualified_request_onchip_memory_s1;
  wire             sgdma_rx_m_write_requests_onchip_memory_s1;
  wire             sgdma_rx_m_write_saved_grant_onchip_memory_s1;
  wire             sgdma_tx_m_read_arbiterlock;
  wire             sgdma_tx_m_read_arbiterlock2;
  wire             sgdma_tx_m_read_continuerequest;
  wire             sgdma_tx_m_read_granted_onchip_memory_s1;
  wire             sgdma_tx_m_read_qualified_request_onchip_memory_s1;
  wire             sgdma_tx_m_read_read_data_valid_onchip_memory_s1;
  reg              sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register;
  wire             sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register_in;
  wire             sgdma_tx_m_read_requests_onchip_memory_s1;
  wire             sgdma_tx_m_read_saved_grant_onchip_memory_s1;
  wire    [ 30: 0] shifted_address_to_onchip_memory_s1_from_cpu_data_master;
  wire    [ 30: 0] shifted_address_to_onchip_memory_s1_from_cpu_instruction_master;
  wire    [ 31: 0] shifted_address_to_onchip_memory_s1_from_sgdma_rx_m_write;
  wire    [ 31: 0] shifted_address_to_onchip_memory_s1_from_sgdma_tx_m_read;
  wire             wait_for_onchip_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~onchip_memory_s1_end_xfer;
    end


  assign onchip_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_onchip_memory_s1 | cpu_instruction_master_qualified_request_onchip_memory_s1 | sgdma_rx_m_write_qualified_request_onchip_memory_s1 | sgdma_tx_m_read_qualified_request_onchip_memory_s1));
  //assign onchip_memory_s1_readdata_from_sa = onchip_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_memory_s1_readdata_from_sa = onchip_memory_s1_readdata;

  assign cpu_data_master_requests_onchip_memory_s1 = ({cpu_data_master_address_to_slave[30 : 19] , 19'b0} == 31'h48080000) & (cpu_data_master_read | cpu_data_master_write);
  //onchip_memory_s1_arb_share_counter set values, which is an e_mux
  assign onchip_memory_s1_arb_share_set_values = 1;

  //onchip_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_memory_s1_non_bursting_master_requests = cpu_data_master_requests_onchip_memory_s1 |
    cpu_instruction_master_requests_onchip_memory_s1 |
    sgdma_rx_m_write_requests_onchip_memory_s1 |
    sgdma_tx_m_read_requests_onchip_memory_s1 |
    cpu_data_master_requests_onchip_memory_s1 |
    cpu_instruction_master_requests_onchip_memory_s1 |
    sgdma_rx_m_write_requests_onchip_memory_s1 |
    sgdma_tx_m_read_requests_onchip_memory_s1 |
    cpu_data_master_requests_onchip_memory_s1 |
    cpu_instruction_master_requests_onchip_memory_s1 |
    sgdma_rx_m_write_requests_onchip_memory_s1 |
    sgdma_tx_m_read_requests_onchip_memory_s1 |
    cpu_data_master_requests_onchip_memory_s1 |
    cpu_instruction_master_requests_onchip_memory_s1 |
    sgdma_rx_m_write_requests_onchip_memory_s1 |
    sgdma_tx_m_read_requests_onchip_memory_s1;

  //onchip_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_memory_s1_any_bursting_master_saved_grant = 0;

  //onchip_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_memory_s1_arb_share_counter_next_value = onchip_memory_s1_firsttransfer ? (onchip_memory_s1_arb_share_set_values - 1) : |onchip_memory_s1_arb_share_counter ? (onchip_memory_s1_arb_share_counter - 1) : 0;

  //onchip_memory_s1_allgrants all slave grants, which is an e_mux
  assign onchip_memory_s1_allgrants = (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector) |
    (|onchip_memory_s1_grant_vector);

  //onchip_memory_s1_end_xfer assignment, which is an e_assign
  assign onchip_memory_s1_end_xfer = ~(onchip_memory_s1_waits_for_read | onchip_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_memory_s1 = onchip_memory_s1_end_xfer & (~onchip_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_memory_s1 & onchip_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_memory_s1 & ~onchip_memory_s1_non_bursting_master_requests);

  //onchip_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory_s1_arb_share_counter <= 0;
      else if (onchip_memory_s1_arb_counter_enable)
          onchip_memory_s1_arb_share_counter <= onchip_memory_s1_arb_share_counter_next_value;
    end


  //onchip_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_memory_s1) | (end_xfer_arb_share_counter_term_onchip_memory_s1 & ~onchip_memory_s1_non_bursting_master_requests))
          onchip_memory_s1_slavearbiterlockenable <= |onchip_memory_s1_arb_share_counter_next_value;
    end


  //cpu/data_master onchip_memory/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = onchip_memory_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //onchip_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_memory_s1_slavearbiterlockenable2 = |onchip_memory_s1_arb_share_counter_next_value;

  //cpu/data_master onchip_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = onchip_memory_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master onchip_memory/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = onchip_memory_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master onchip_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = onchip_memory_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted onchip_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1 <= cpu_instruction_master_saved_grant_onchip_memory_s1 ? 1 : (onchip_memory_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_onchip_memory_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = (last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1 & cpu_instruction_master_requests_onchip_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1 & cpu_instruction_master_requests_onchip_memory_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_onchip_memory_s1 & cpu_instruction_master_requests_onchip_memory_s1);

  //onchip_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_memory_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    sgdma_rx_m_write_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_m_write_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write onchip_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock = onchip_memory_s1_slavearbiterlockenable & sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write onchip_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock2 = onchip_memory_s1_slavearbiterlockenable2 & sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write granted onchip_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1 <= sgdma_rx_m_write_saved_grant_onchip_memory_s1 ? 1 : (onchip_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_m_write_requests_onchip_memory_s1) ? 0 : last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1;
    end


  //sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_m_write_continuerequest = (last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1 & sgdma_rx_m_write_requests_onchip_memory_s1) |
    (last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1 & sgdma_rx_m_write_requests_onchip_memory_s1) |
    (last_cycle_sgdma_rx_m_write_granted_slave_onchip_memory_s1 & sgdma_rx_m_write_requests_onchip_memory_s1);

  //sgdma_tx/m_read onchip_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock = onchip_memory_s1_slavearbiterlockenable & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read onchip_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock2 = onchip_memory_s1_slavearbiterlockenable2 & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read granted onchip_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1 <= sgdma_tx_m_read_saved_grant_onchip_memory_s1 ? 1 : (onchip_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_m_read_requests_onchip_memory_s1) ? 0 : last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1;
    end


  //sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_m_read_continuerequest = (last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1 & sgdma_tx_m_read_requests_onchip_memory_s1) |
    (last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1 & sgdma_tx_m_read_requests_onchip_memory_s1) |
    (last_cycle_sgdma_tx_m_read_granted_slave_onchip_memory_s1 & sgdma_tx_m_read_requests_onchip_memory_s1);

  assign cpu_data_master_qualified_request_onchip_memory_s1 = cpu_data_master_requests_onchip_memory_s1 & ~((cpu_data_master_read & ((1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))) | cpu_instruction_master_arbiterlock | sgdma_rx_m_write_arbiterlock | sgdma_tx_m_read_arbiterlock);
  //cpu_data_master_read_data_valid_onchip_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_data_master_read_data_valid_onchip_memory_s1_shift_register_in = cpu_data_master_granted_onchip_memory_s1 & cpu_data_master_read & ~onchip_memory_s1_waits_for_read;

  //shift register p1 cpu_data_master_read_data_valid_onchip_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_data_master_read_data_valid_onchip_memory_s1_shift_register = {cpu_data_master_read_data_valid_onchip_memory_s1_shift_register, cpu_data_master_read_data_valid_onchip_memory_s1_shift_register_in};

  //cpu_data_master_read_data_valid_onchip_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_data_valid_onchip_memory_s1_shift_register <= 0;
      else 
        cpu_data_master_read_data_valid_onchip_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_onchip_memory_s1_shift_register;
    end


  //local readdatavalid cpu_data_master_read_data_valid_onchip_memory_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_onchip_memory_s1 = cpu_data_master_read_data_valid_onchip_memory_s1_shift_register;

  //onchip_memory_s1_writedata mux, which is an e_mux
  assign onchip_memory_s1_writedata = (cpu_data_master_granted_onchip_memory_s1)? cpu_data_master_writedata :
    sgdma_rx_m_write_writedata;

  //mux onchip_memory_s1_clken, which is an e_mux
  assign onchip_memory_s1_clken = 1'b1;

  assign cpu_instruction_master_requests_onchip_memory_s1 = (({cpu_instruction_master_address_to_slave[30 : 19] , 19'b0} == 31'h48080000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted onchip_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_onchip_memory_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_onchip_memory_s1 <= cpu_data_master_saved_grant_onchip_memory_s1 ? 1 : (onchip_memory_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_onchip_memory_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_onchip_memory_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = (last_cycle_cpu_data_master_granted_slave_onchip_memory_s1 & cpu_data_master_requests_onchip_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_onchip_memory_s1 & cpu_data_master_requests_onchip_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_onchip_memory_s1 & cpu_data_master_requests_onchip_memory_s1);

  assign cpu_instruction_master_qualified_request_onchip_memory_s1 = cpu_instruction_master_requests_onchip_memory_s1 & ~((cpu_instruction_master_read & ((1 < cpu_instruction_master_latency_counter))) | cpu_data_master_arbiterlock | sgdma_rx_m_write_arbiterlock | sgdma_tx_m_read_arbiterlock);
  //cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in = cpu_instruction_master_granted_onchip_memory_s1 & cpu_instruction_master_read & ~onchip_memory_s1_waits_for_read;

  //shift register p1 cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register = {cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register, cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in};

  //cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register <= 0;
      else 
        cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register <= p1_cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register;
    end


  //local readdatavalid cpu_instruction_master_read_data_valid_onchip_memory_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_onchip_memory_s1 = cpu_instruction_master_read_data_valid_onchip_memory_s1_shift_register;

  assign sgdma_rx_m_write_requests_onchip_memory_s1 = (({sgdma_rx_m_write_address_to_slave[31 : 19] , 19'b0} == 32'h48080000) & (sgdma_rx_m_write_write)) & sgdma_rx_m_write_write;
  assign sgdma_rx_m_write_qualified_request_onchip_memory_s1 = sgdma_rx_m_write_requests_onchip_memory_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_tx_m_read_arbiterlock);
  assign sgdma_tx_m_read_requests_onchip_memory_s1 = (({sgdma_tx_m_read_address_to_slave[31 : 19] , 19'b0} == 32'h48080000) & (sgdma_tx_m_read_read)) & sgdma_tx_m_read_read;
  assign sgdma_tx_m_read_qualified_request_onchip_memory_s1 = sgdma_tx_m_read_requests_onchip_memory_s1 & ~((sgdma_tx_m_read_read & ((1 < sgdma_tx_m_read_latency_counter))) | cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_m_write_arbiterlock);
  //sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register_in = sgdma_tx_m_read_granted_onchip_memory_s1 & sgdma_tx_m_read_read & ~onchip_memory_s1_waits_for_read;

  //shift register p1 sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register = {sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register, sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register_in};

  //sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register <= 0;
      else 
        sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register <= p1_sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register;
    end


  //local readdatavalid sgdma_tx_m_read_read_data_valid_onchip_memory_s1, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_onchip_memory_s1 = sgdma_tx_m_read_read_data_valid_onchip_memory_s1_shift_register;

  //allow new arb cycle for onchip_memory/s1, which is an e_assign
  assign onchip_memory_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock & ~sgdma_rx_m_write_arbiterlock & ~sgdma_tx_m_read_arbiterlock;

  //sgdma_tx/m_read assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  assign onchip_memory_s1_master_qreq_vector[0] = sgdma_tx_m_read_qualified_request_onchip_memory_s1;

  //sgdma_tx/m_read grant onchip_memory/s1, which is an e_assign
  assign sgdma_tx_m_read_granted_onchip_memory_s1 = onchip_memory_s1_grant_vector[0];

  //sgdma_tx/m_read saved-grant onchip_memory/s1, which is an e_assign
  assign sgdma_tx_m_read_saved_grant_onchip_memory_s1 = onchip_memory_s1_arb_winner[0] && sgdma_tx_m_read_requests_onchip_memory_s1;

  //sgdma_rx/m_write assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  assign onchip_memory_s1_master_qreq_vector[1] = sgdma_rx_m_write_qualified_request_onchip_memory_s1;

  //sgdma_rx/m_write grant onchip_memory/s1, which is an e_assign
  assign sgdma_rx_m_write_granted_onchip_memory_s1 = onchip_memory_s1_grant_vector[1];

  //sgdma_rx/m_write saved-grant onchip_memory/s1, which is an e_assign
  assign sgdma_rx_m_write_saved_grant_onchip_memory_s1 = onchip_memory_s1_arb_winner[1] && sgdma_rx_m_write_requests_onchip_memory_s1;

  //cpu/instruction_master assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  assign onchip_memory_s1_master_qreq_vector[2] = cpu_instruction_master_qualified_request_onchip_memory_s1;

  //cpu/instruction_master grant onchip_memory/s1, which is an e_assign
  assign cpu_instruction_master_granted_onchip_memory_s1 = onchip_memory_s1_grant_vector[2];

  //cpu/instruction_master saved-grant onchip_memory/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_onchip_memory_s1 = onchip_memory_s1_arb_winner[2] && cpu_instruction_master_requests_onchip_memory_s1;

  //cpu/data_master assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  assign onchip_memory_s1_master_qreq_vector[3] = cpu_data_master_qualified_request_onchip_memory_s1;

  //cpu/data_master grant onchip_memory/s1, which is an e_assign
  assign cpu_data_master_granted_onchip_memory_s1 = onchip_memory_s1_grant_vector[3];

  //cpu/data_master saved-grant onchip_memory/s1, which is an e_assign
  assign cpu_data_master_saved_grant_onchip_memory_s1 = onchip_memory_s1_arb_winner[3] && cpu_data_master_requests_onchip_memory_s1;

  //onchip_memory/s1 chosen-master double-vector, which is an e_assign
  assign onchip_memory_s1_chosen_master_double_vector = {onchip_memory_s1_master_qreq_vector, onchip_memory_s1_master_qreq_vector} & ({~onchip_memory_s1_master_qreq_vector, ~onchip_memory_s1_master_qreq_vector} + onchip_memory_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_memory_s1_arb_winner = (onchip_memory_s1_allow_new_arb_cycle & | onchip_memory_s1_grant_vector) ? onchip_memory_s1_grant_vector : onchip_memory_s1_saved_chosen_master_vector;

  //saved onchip_memory_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory_s1_saved_chosen_master_vector <= 0;
      else if (onchip_memory_s1_allow_new_arb_cycle)
          onchip_memory_s1_saved_chosen_master_vector <= |onchip_memory_s1_grant_vector ? onchip_memory_s1_grant_vector : onchip_memory_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_memory_s1_grant_vector = {(onchip_memory_s1_chosen_master_double_vector[3] | onchip_memory_s1_chosen_master_double_vector[7]),
    (onchip_memory_s1_chosen_master_double_vector[2] | onchip_memory_s1_chosen_master_double_vector[6]),
    (onchip_memory_s1_chosen_master_double_vector[1] | onchip_memory_s1_chosen_master_double_vector[5]),
    (onchip_memory_s1_chosen_master_double_vector[0] | onchip_memory_s1_chosen_master_double_vector[4])};

  //onchip_memory/s1 chosen master rotated left, which is an e_assign
  assign onchip_memory_s1_chosen_master_rot_left = (onchip_memory_s1_arb_winner << 1) ? (onchip_memory_s1_arb_winner << 1) : 1;

  //onchip_memory/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory_s1_arb_addend <= 1;
      else if (|onchip_memory_s1_grant_vector)
          onchip_memory_s1_arb_addend <= onchip_memory_s1_end_xfer? onchip_memory_s1_chosen_master_rot_left : onchip_memory_s1_grant_vector;
    end


  assign onchip_memory_s1_chipselect = cpu_data_master_granted_onchip_memory_s1 | cpu_instruction_master_granted_onchip_memory_s1 | sgdma_rx_m_write_granted_onchip_memory_s1 | sgdma_tx_m_read_granted_onchip_memory_s1;
  //onchip_memory_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_memory_s1_firsttransfer = onchip_memory_s1_begins_xfer ? onchip_memory_s1_unreg_firsttransfer : onchip_memory_s1_reg_firsttransfer;

  //onchip_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_memory_s1_unreg_firsttransfer = ~(onchip_memory_s1_slavearbiterlockenable & onchip_memory_s1_any_continuerequest);

  //onchip_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_memory_s1_begins_xfer)
          onchip_memory_s1_reg_firsttransfer <= onchip_memory_s1_unreg_firsttransfer;
    end


  //onchip_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_memory_s1_beginbursttransfer_internal = onchip_memory_s1_begins_xfer;

  //onchip_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_memory_s1_arbitration_holdoff_internal = onchip_memory_s1_begins_xfer & onchip_memory_s1_firsttransfer;

  //onchip_memory_s1_write assignment, which is an e_mux
  assign onchip_memory_s1_write = (cpu_data_master_granted_onchip_memory_s1 & cpu_data_master_write) | (sgdma_rx_m_write_granted_onchip_memory_s1 & sgdma_rx_m_write_write);

  assign shifted_address_to_onchip_memory_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //onchip_memory_s1_address mux, which is an e_mux
  assign onchip_memory_s1_address = (cpu_data_master_granted_onchip_memory_s1)? (shifted_address_to_onchip_memory_s1_from_cpu_data_master >> 2) :
    (cpu_instruction_master_granted_onchip_memory_s1)? (shifted_address_to_onchip_memory_s1_from_cpu_instruction_master >> 2) :
    (sgdma_rx_m_write_granted_onchip_memory_s1)? (shifted_address_to_onchip_memory_s1_from_sgdma_rx_m_write >> 2) :
    (shifted_address_to_onchip_memory_s1_from_sgdma_tx_m_read >> 2);

  assign shifted_address_to_onchip_memory_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory_s1_from_sgdma_rx_m_write = sgdma_rx_m_write_address_to_slave;
  assign shifted_address_to_onchip_memory_s1_from_sgdma_tx_m_read = sgdma_tx_m_read_address_to_slave;
  //d1_onchip_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_memory_s1_end_xfer <= 1;
      else 
        d1_onchip_memory_s1_end_xfer <= onchip_memory_s1_end_xfer;
    end


  //onchip_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_memory_s1_waits_for_read = onchip_memory_s1_in_a_read_cycle & 0;

  //onchip_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_memory_s1_in_a_read_cycle = (cpu_data_master_granted_onchip_memory_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_onchip_memory_s1 & cpu_instruction_master_read) | (sgdma_tx_m_read_granted_onchip_memory_s1 & sgdma_tx_m_read_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_memory_s1_in_a_read_cycle;

  //onchip_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_memory_s1_waits_for_write = onchip_memory_s1_in_a_write_cycle & 0;

  //onchip_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_memory_s1_in_a_write_cycle = (cpu_data_master_granted_onchip_memory_s1 & cpu_data_master_write) | (sgdma_rx_m_write_granted_onchip_memory_s1 & sgdma_rx_m_write_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_memory_s1_in_a_write_cycle;

  assign wait_for_onchip_memory_s1_counter = 0;
  //onchip_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_memory_s1_byteenable = (cpu_data_master_granted_onchip_memory_s1)? cpu_data_master_byteenable :
    (sgdma_rx_m_write_granted_onchip_memory_s1)? sgdma_rx_m_write_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_onchip_memory_s1 + cpu_instruction_master_granted_onchip_memory_s1 + sgdma_rx_m_write_granted_onchip_memory_s1 + sgdma_tx_m_read_granted_onchip_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_onchip_memory_s1 + cpu_instruction_master_saved_grant_onchip_memory_s1 + sgdma_rx_m_write_saved_grant_onchip_memory_s1 + sgdma_tx_m_read_saved_grant_onchip_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module packet_memory_s1_arbitrator (
                                     // inputs:
                                      clk,
                                      cpu_data_master_address_to_slave,
                                      cpu_data_master_byteenable,
                                      cpu_data_master_latency_counter,
                                      cpu_data_master_read,
                                      cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                      cpu_data_master_write,
                                      cpu_data_master_writedata,
                                      packet_memory_s1_readdata,
                                      reset_n,

                                     // outputs:
                                      cpu_data_master_granted_packet_memory_s1,
                                      cpu_data_master_qualified_request_packet_memory_s1,
                                      cpu_data_master_read_data_valid_packet_memory_s1,
                                      cpu_data_master_requests_packet_memory_s1,
                                      d1_packet_memory_s1_end_xfer,
                                      packet_memory_s1_address,
                                      packet_memory_s1_byteenable,
                                      packet_memory_s1_chipselect,
                                      packet_memory_s1_clken,
                                      packet_memory_s1_readdata_from_sa,
                                      packet_memory_s1_write,
                                      packet_memory_s1_writedata
                                   )
;

  output           cpu_data_master_granted_packet_memory_s1;
  output           cpu_data_master_qualified_request_packet_memory_s1;
  output           cpu_data_master_read_data_valid_packet_memory_s1;
  output           cpu_data_master_requests_packet_memory_s1;
  output           d1_packet_memory_s1_end_xfer;
  output  [ 13: 0] packet_memory_s1_address;
  output  [  3: 0] packet_memory_s1_byteenable;
  output           packet_memory_s1_chipselect;
  output           packet_memory_s1_clken;
  output  [ 31: 0] packet_memory_s1_readdata_from_sa;
  output           packet_memory_s1_write;
  output  [ 31: 0] packet_memory_s1_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] packet_memory_s1_readdata;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_packet_memory_s1;
  wire             cpu_data_master_qualified_request_packet_memory_s1;
  wire             cpu_data_master_read_data_valid_packet_memory_s1;
  reg              cpu_data_master_read_data_valid_packet_memory_s1_shift_register;
  wire             cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in;
  wire             cpu_data_master_requests_packet_memory_s1;
  wire             cpu_data_master_saved_grant_packet_memory_s1;
  reg              d1_packet_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_packet_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register;
  wire    [ 13: 0] packet_memory_s1_address;
  wire             packet_memory_s1_allgrants;
  wire             packet_memory_s1_allow_new_arb_cycle;
  wire             packet_memory_s1_any_bursting_master_saved_grant;
  wire             packet_memory_s1_any_continuerequest;
  wire             packet_memory_s1_arb_counter_enable;
  reg     [  1: 0] packet_memory_s1_arb_share_counter;
  wire    [  1: 0] packet_memory_s1_arb_share_counter_next_value;
  wire    [  1: 0] packet_memory_s1_arb_share_set_values;
  wire             packet_memory_s1_beginbursttransfer_internal;
  wire             packet_memory_s1_begins_xfer;
  wire    [  3: 0] packet_memory_s1_byteenable;
  wire             packet_memory_s1_chipselect;
  wire             packet_memory_s1_clken;
  wire             packet_memory_s1_end_xfer;
  wire             packet_memory_s1_firsttransfer;
  wire             packet_memory_s1_grant_vector;
  wire             packet_memory_s1_in_a_read_cycle;
  wire             packet_memory_s1_in_a_write_cycle;
  wire             packet_memory_s1_master_qreq_vector;
  wire             packet_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] packet_memory_s1_readdata_from_sa;
  reg              packet_memory_s1_reg_firsttransfer;
  reg              packet_memory_s1_slavearbiterlockenable;
  wire             packet_memory_s1_slavearbiterlockenable2;
  wire             packet_memory_s1_unreg_firsttransfer;
  wire             packet_memory_s1_waits_for_read;
  wire             packet_memory_s1_waits_for_write;
  wire             packet_memory_s1_write;
  wire    [ 31: 0] packet_memory_s1_writedata;
  wire    [ 30: 0] shifted_address_to_packet_memory_s1_from_cpu_data_master;
  wire             wait_for_packet_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~packet_memory_s1_end_xfer;
    end


  assign packet_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_packet_memory_s1));
  //assign packet_memory_s1_readdata_from_sa = packet_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign packet_memory_s1_readdata_from_sa = packet_memory_s1_readdata;

  assign cpu_data_master_requests_packet_memory_s1 = ({cpu_data_master_address_to_slave[30 : 16] , 16'b0} == 31'h48100000) & (cpu_data_master_read | cpu_data_master_write);
  //packet_memory_s1_arb_share_counter set values, which is an e_mux
  assign packet_memory_s1_arb_share_set_values = 1;

  //packet_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign packet_memory_s1_non_bursting_master_requests = cpu_data_master_requests_packet_memory_s1;

  //packet_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign packet_memory_s1_any_bursting_master_saved_grant = 0;

  //packet_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign packet_memory_s1_arb_share_counter_next_value = packet_memory_s1_firsttransfer ? (packet_memory_s1_arb_share_set_values - 1) : |packet_memory_s1_arb_share_counter ? (packet_memory_s1_arb_share_counter - 1) : 0;

  //packet_memory_s1_allgrants all slave grants, which is an e_mux
  assign packet_memory_s1_allgrants = |packet_memory_s1_grant_vector;

  //packet_memory_s1_end_xfer assignment, which is an e_assign
  assign packet_memory_s1_end_xfer = ~(packet_memory_s1_waits_for_read | packet_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_packet_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_packet_memory_s1 = packet_memory_s1_end_xfer & (~packet_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //packet_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign packet_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_packet_memory_s1 & packet_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_packet_memory_s1 & ~packet_memory_s1_non_bursting_master_requests);

  //packet_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s1_arb_share_counter <= 0;
      else if (packet_memory_s1_arb_counter_enable)
          packet_memory_s1_arb_share_counter <= packet_memory_s1_arb_share_counter_next_value;
    end


  //packet_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s1_slavearbiterlockenable <= 0;
      else if ((|packet_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_packet_memory_s1) | (end_xfer_arb_share_counter_term_packet_memory_s1 & ~packet_memory_s1_non_bursting_master_requests))
          packet_memory_s1_slavearbiterlockenable <= |packet_memory_s1_arb_share_counter_next_value;
    end


  //cpu/data_master packet_memory/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = packet_memory_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //packet_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign packet_memory_s1_slavearbiterlockenable2 = |packet_memory_s1_arb_share_counter_next_value;

  //cpu/data_master packet_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = packet_memory_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //packet_memory_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign packet_memory_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_packet_memory_s1 = cpu_data_master_requests_packet_memory_s1 & ~((cpu_data_master_read & ((1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in = cpu_data_master_granted_packet_memory_s1 & cpu_data_master_read & ~packet_memory_s1_waits_for_read;

  //shift register p1 cpu_data_master_read_data_valid_packet_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register = {cpu_data_master_read_data_valid_packet_memory_s1_shift_register, cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in};

  //cpu_data_master_read_data_valid_packet_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_data_valid_packet_memory_s1_shift_register <= 0;
      else 
        cpu_data_master_read_data_valid_packet_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register;
    end


  //local readdatavalid cpu_data_master_read_data_valid_packet_memory_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_packet_memory_s1 = cpu_data_master_read_data_valid_packet_memory_s1_shift_register;

  //packet_memory_s1_writedata mux, which is an e_mux
  assign packet_memory_s1_writedata = cpu_data_master_writedata;

  //mux packet_memory_s1_clken, which is an e_mux
  assign packet_memory_s1_clken = 1'b1;

  //master is always granted when requested
  assign cpu_data_master_granted_packet_memory_s1 = cpu_data_master_qualified_request_packet_memory_s1;

  //cpu/data_master saved-grant packet_memory/s1, which is an e_assign
  assign cpu_data_master_saved_grant_packet_memory_s1 = cpu_data_master_requests_packet_memory_s1;

  //allow new arb cycle for packet_memory/s1, which is an e_assign
  assign packet_memory_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign packet_memory_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign packet_memory_s1_master_qreq_vector = 1;

  assign packet_memory_s1_chipselect = cpu_data_master_granted_packet_memory_s1;
  //packet_memory_s1_firsttransfer first transaction, which is an e_assign
  assign packet_memory_s1_firsttransfer = packet_memory_s1_begins_xfer ? packet_memory_s1_unreg_firsttransfer : packet_memory_s1_reg_firsttransfer;

  //packet_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign packet_memory_s1_unreg_firsttransfer = ~(packet_memory_s1_slavearbiterlockenable & packet_memory_s1_any_continuerequest);

  //packet_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s1_reg_firsttransfer <= 1'b1;
      else if (packet_memory_s1_begins_xfer)
          packet_memory_s1_reg_firsttransfer <= packet_memory_s1_unreg_firsttransfer;
    end


  //packet_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign packet_memory_s1_beginbursttransfer_internal = packet_memory_s1_begins_xfer;

  //packet_memory_s1_write assignment, which is an e_mux
  assign packet_memory_s1_write = cpu_data_master_granted_packet_memory_s1 & cpu_data_master_write;

  assign shifted_address_to_packet_memory_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //packet_memory_s1_address mux, which is an e_mux
  assign packet_memory_s1_address = shifted_address_to_packet_memory_s1_from_cpu_data_master >> 2;

  //d1_packet_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_packet_memory_s1_end_xfer <= 1;
      else 
        d1_packet_memory_s1_end_xfer <= packet_memory_s1_end_xfer;
    end


  //packet_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign packet_memory_s1_waits_for_read = packet_memory_s1_in_a_read_cycle & 0;

  //packet_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign packet_memory_s1_in_a_read_cycle = cpu_data_master_granted_packet_memory_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = packet_memory_s1_in_a_read_cycle;

  //packet_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign packet_memory_s1_waits_for_write = packet_memory_s1_in_a_write_cycle & 0;

  //packet_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign packet_memory_s1_in_a_write_cycle = cpu_data_master_granted_packet_memory_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = packet_memory_s1_in_a_write_cycle;

  assign wait_for_packet_memory_s1_counter = 0;
  //packet_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign packet_memory_s1_byteenable = (cpu_data_master_granted_packet_memory_s1)? cpu_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //packet_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module packet_memory_s2_arbitrator (
                                     // inputs:
                                      clk,
                                      packet_memory_s2_readdata,
                                      reset_n,
                                      sgdma_rx_m_write_address_to_slave,
                                      sgdma_rx_m_write_byteenable,
                                      sgdma_rx_m_write_write,
                                      sgdma_rx_m_write_writedata,
                                      sgdma_tx_m_read_address_to_slave,
                                      sgdma_tx_m_read_latency_counter,
                                      sgdma_tx_m_read_read,

                                     // outputs:
                                      d1_packet_memory_s2_end_xfer,
                                      packet_memory_s2_address,
                                      packet_memory_s2_byteenable,
                                      packet_memory_s2_chipselect,
                                      packet_memory_s2_clken,
                                      packet_memory_s2_readdata_from_sa,
                                      packet_memory_s2_write,
                                      packet_memory_s2_writedata,
                                      sgdma_rx_m_write_granted_packet_memory_s2,
                                      sgdma_rx_m_write_qualified_request_packet_memory_s2,
                                      sgdma_rx_m_write_requests_packet_memory_s2,
                                      sgdma_tx_m_read_granted_packet_memory_s2,
                                      sgdma_tx_m_read_qualified_request_packet_memory_s2,
                                      sgdma_tx_m_read_read_data_valid_packet_memory_s2,
                                      sgdma_tx_m_read_requests_packet_memory_s2
                                   )
;

  output           d1_packet_memory_s2_end_xfer;
  output  [ 13: 0] packet_memory_s2_address;
  output  [  3: 0] packet_memory_s2_byteenable;
  output           packet_memory_s2_chipselect;
  output           packet_memory_s2_clken;
  output  [ 31: 0] packet_memory_s2_readdata_from_sa;
  output           packet_memory_s2_write;
  output  [ 31: 0] packet_memory_s2_writedata;
  output           sgdma_rx_m_write_granted_packet_memory_s2;
  output           sgdma_rx_m_write_qualified_request_packet_memory_s2;
  output           sgdma_rx_m_write_requests_packet_memory_s2;
  output           sgdma_tx_m_read_granted_packet_memory_s2;
  output           sgdma_tx_m_read_qualified_request_packet_memory_s2;
  output           sgdma_tx_m_read_read_data_valid_packet_memory_s2;
  output           sgdma_tx_m_read_requests_packet_memory_s2;
  input            clk;
  input   [ 31: 0] packet_memory_s2_readdata;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address_to_slave;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;
  input   [ 31: 0] sgdma_tx_m_read_address_to_slave;
  input            sgdma_tx_m_read_latency_counter;
  input            sgdma_tx_m_read_read;

  reg              d1_packet_memory_s2_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_packet_memory_s2;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2;
  reg              last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2;
  wire             p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;
  wire    [ 13: 0] packet_memory_s2_address;
  wire             packet_memory_s2_allgrants;
  wire             packet_memory_s2_allow_new_arb_cycle;
  wire             packet_memory_s2_any_bursting_master_saved_grant;
  wire             packet_memory_s2_any_continuerequest;
  reg     [  1: 0] packet_memory_s2_arb_addend;
  wire             packet_memory_s2_arb_counter_enable;
  reg              packet_memory_s2_arb_share_counter;
  wire             packet_memory_s2_arb_share_counter_next_value;
  wire             packet_memory_s2_arb_share_set_values;
  wire    [  1: 0] packet_memory_s2_arb_winner;
  wire             packet_memory_s2_arbitration_holdoff_internal;
  wire             packet_memory_s2_beginbursttransfer_internal;
  wire             packet_memory_s2_begins_xfer;
  wire    [  3: 0] packet_memory_s2_byteenable;
  wire             packet_memory_s2_chipselect;
  wire    [  3: 0] packet_memory_s2_chosen_master_double_vector;
  wire    [  1: 0] packet_memory_s2_chosen_master_rot_left;
  wire             packet_memory_s2_clken;
  wire             packet_memory_s2_end_xfer;
  wire             packet_memory_s2_firsttransfer;
  wire    [  1: 0] packet_memory_s2_grant_vector;
  wire             packet_memory_s2_in_a_read_cycle;
  wire             packet_memory_s2_in_a_write_cycle;
  wire    [  1: 0] packet_memory_s2_master_qreq_vector;
  wire             packet_memory_s2_non_bursting_master_requests;
  wire    [ 31: 0] packet_memory_s2_readdata_from_sa;
  reg              packet_memory_s2_reg_firsttransfer;
  reg     [  1: 0] packet_memory_s2_saved_chosen_master_vector;
  reg              packet_memory_s2_slavearbiterlockenable;
  wire             packet_memory_s2_slavearbiterlockenable2;
  wire             packet_memory_s2_unreg_firsttransfer;
  wire             packet_memory_s2_waits_for_read;
  wire             packet_memory_s2_waits_for_write;
  wire             packet_memory_s2_write;
  wire    [ 31: 0] packet_memory_s2_writedata;
  wire             sgdma_rx_m_write_arbiterlock;
  wire             sgdma_rx_m_write_arbiterlock2;
  wire             sgdma_rx_m_write_continuerequest;
  wire             sgdma_rx_m_write_granted_packet_memory_s2;
  wire             sgdma_rx_m_write_qualified_request_packet_memory_s2;
  wire             sgdma_rx_m_write_requests_packet_memory_s2;
  wire             sgdma_rx_m_write_saved_grant_packet_memory_s2;
  wire             sgdma_tx_m_read_arbiterlock;
  wire             sgdma_tx_m_read_arbiterlock2;
  wire             sgdma_tx_m_read_continuerequest;
  wire             sgdma_tx_m_read_granted_packet_memory_s2;
  wire             sgdma_tx_m_read_qualified_request_packet_memory_s2;
  wire             sgdma_tx_m_read_read_data_valid_packet_memory_s2;
  reg              sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;
  wire             sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in;
  wire             sgdma_tx_m_read_requests_packet_memory_s2;
  wire             sgdma_tx_m_read_saved_grant_packet_memory_s2;
  wire    [ 31: 0] shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write;
  wire    [ 31: 0] shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read;
  wire             wait_for_packet_memory_s2_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~packet_memory_s2_end_xfer;
    end


  assign packet_memory_s2_begins_xfer = ~d1_reasons_to_wait & ((sgdma_rx_m_write_qualified_request_packet_memory_s2 | sgdma_tx_m_read_qualified_request_packet_memory_s2));
  //assign packet_memory_s2_readdata_from_sa = packet_memory_s2_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign packet_memory_s2_readdata_from_sa = packet_memory_s2_readdata;

  assign sgdma_rx_m_write_requests_packet_memory_s2 = (({sgdma_rx_m_write_address_to_slave[31 : 16] , 16'b0} == 32'h48100000) & (sgdma_rx_m_write_write)) & sgdma_rx_m_write_write;
  //packet_memory_s2_arb_share_counter set values, which is an e_mux
  assign packet_memory_s2_arb_share_set_values = 1;

  //packet_memory_s2_non_bursting_master_requests mux, which is an e_mux
  assign packet_memory_s2_non_bursting_master_requests = sgdma_rx_m_write_requests_packet_memory_s2 |
    sgdma_tx_m_read_requests_packet_memory_s2 |
    sgdma_rx_m_write_requests_packet_memory_s2 |
    sgdma_tx_m_read_requests_packet_memory_s2;

  //packet_memory_s2_any_bursting_master_saved_grant mux, which is an e_mux
  assign packet_memory_s2_any_bursting_master_saved_grant = 0;

  //packet_memory_s2_arb_share_counter_next_value assignment, which is an e_assign
  assign packet_memory_s2_arb_share_counter_next_value = packet_memory_s2_firsttransfer ? (packet_memory_s2_arb_share_set_values - 1) : |packet_memory_s2_arb_share_counter ? (packet_memory_s2_arb_share_counter - 1) : 0;

  //packet_memory_s2_allgrants all slave grants, which is an e_mux
  assign packet_memory_s2_allgrants = (|packet_memory_s2_grant_vector) |
    (|packet_memory_s2_grant_vector) |
    (|packet_memory_s2_grant_vector) |
    (|packet_memory_s2_grant_vector);

  //packet_memory_s2_end_xfer assignment, which is an e_assign
  assign packet_memory_s2_end_xfer = ~(packet_memory_s2_waits_for_read | packet_memory_s2_waits_for_write);

  //end_xfer_arb_share_counter_term_packet_memory_s2 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_packet_memory_s2 = packet_memory_s2_end_xfer & (~packet_memory_s2_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //packet_memory_s2_arb_share_counter arbitration counter enable, which is an e_assign
  assign packet_memory_s2_arb_counter_enable = (end_xfer_arb_share_counter_term_packet_memory_s2 & packet_memory_s2_allgrants) | (end_xfer_arb_share_counter_term_packet_memory_s2 & ~packet_memory_s2_non_bursting_master_requests);

  //packet_memory_s2_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s2_arb_share_counter <= 0;
      else if (packet_memory_s2_arb_counter_enable)
          packet_memory_s2_arb_share_counter <= packet_memory_s2_arb_share_counter_next_value;
    end


  //packet_memory_s2_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s2_slavearbiterlockenable <= 0;
      else if ((|packet_memory_s2_master_qreq_vector & end_xfer_arb_share_counter_term_packet_memory_s2) | (end_xfer_arb_share_counter_term_packet_memory_s2 & ~packet_memory_s2_non_bursting_master_requests))
          packet_memory_s2_slavearbiterlockenable <= |packet_memory_s2_arb_share_counter_next_value;
    end


  //sgdma_rx/m_write packet_memory/s2 arbiterlock, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock = packet_memory_s2_slavearbiterlockenable & sgdma_rx_m_write_continuerequest;

  //packet_memory_s2_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign packet_memory_s2_slavearbiterlockenable2 = |packet_memory_s2_arb_share_counter_next_value;

  //sgdma_rx/m_write packet_memory/s2 arbiterlock2, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock2 = packet_memory_s2_slavearbiterlockenable2 & sgdma_rx_m_write_continuerequest;

  //sgdma_tx/m_read packet_memory/s2 arbiterlock, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock = packet_memory_s2_slavearbiterlockenable & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read packet_memory/s2 arbiterlock2, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock2 = packet_memory_s2_slavearbiterlockenable2 & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read granted packet_memory/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 <= 0;
      else 
        last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 <= sgdma_tx_m_read_saved_grant_packet_memory_s2 ? 1 : (packet_memory_s2_arbitration_holdoff_internal | ~sgdma_tx_m_read_requests_packet_memory_s2) ? 0 : last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2;
    end


  //sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_m_read_continuerequest = last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 & sgdma_tx_m_read_requests_packet_memory_s2;

  //packet_memory_s2_any_continuerequest at least one master continues requesting, which is an e_mux
  assign packet_memory_s2_any_continuerequest = sgdma_tx_m_read_continuerequest |
    sgdma_rx_m_write_continuerequest;

  assign sgdma_rx_m_write_qualified_request_packet_memory_s2 = sgdma_rx_m_write_requests_packet_memory_s2 & ~(sgdma_tx_m_read_arbiterlock);
  //packet_memory_s2_writedata mux, which is an e_mux
  assign packet_memory_s2_writedata = sgdma_rx_m_write_writedata;

  //mux packet_memory_s2_clken, which is an e_mux
  assign packet_memory_s2_clken = 1'b1;

  assign sgdma_tx_m_read_requests_packet_memory_s2 = (({sgdma_tx_m_read_address_to_slave[31 : 16] , 16'b0} == 32'h48100000) & (sgdma_tx_m_read_read)) & sgdma_tx_m_read_read;
  //sgdma_rx/m_write granted packet_memory/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 <= 0;
      else 
        last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 <= sgdma_rx_m_write_saved_grant_packet_memory_s2 ? 1 : (packet_memory_s2_arbitration_holdoff_internal | ~sgdma_rx_m_write_requests_packet_memory_s2) ? 0 : last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2;
    end


  //sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_m_write_continuerequest = last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 & sgdma_rx_m_write_requests_packet_memory_s2;

  assign sgdma_tx_m_read_qualified_request_packet_memory_s2 = sgdma_tx_m_read_requests_packet_memory_s2 & ~((sgdma_tx_m_read_read & ((1 < sgdma_tx_m_read_latency_counter))) | sgdma_rx_m_write_arbiterlock);
  //sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in = sgdma_tx_m_read_granted_packet_memory_s2 & sgdma_tx_m_read_read & ~packet_memory_s2_waits_for_read;

  //shift register p1 sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register = {sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register, sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in};

  //sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register <= 0;
      else 
        sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register <= p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;
    end


  //local readdatavalid sgdma_tx_m_read_read_data_valid_packet_memory_s2, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_packet_memory_s2 = sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;

  //allow new arb cycle for packet_memory/s2, which is an e_assign
  assign packet_memory_s2_allow_new_arb_cycle = ~sgdma_rx_m_write_arbiterlock & ~sgdma_tx_m_read_arbiterlock;

  //sgdma_tx/m_read assignment into master qualified-requests vector for packet_memory/s2, which is an e_assign
  assign packet_memory_s2_master_qreq_vector[0] = sgdma_tx_m_read_qualified_request_packet_memory_s2;

  //sgdma_tx/m_read grant packet_memory/s2, which is an e_assign
  assign sgdma_tx_m_read_granted_packet_memory_s2 = packet_memory_s2_grant_vector[0];

  //sgdma_tx/m_read saved-grant packet_memory/s2, which is an e_assign
  assign sgdma_tx_m_read_saved_grant_packet_memory_s2 = packet_memory_s2_arb_winner[0] && sgdma_tx_m_read_requests_packet_memory_s2;

  //sgdma_rx/m_write assignment into master qualified-requests vector for packet_memory/s2, which is an e_assign
  assign packet_memory_s2_master_qreq_vector[1] = sgdma_rx_m_write_qualified_request_packet_memory_s2;

  //sgdma_rx/m_write grant packet_memory/s2, which is an e_assign
  assign sgdma_rx_m_write_granted_packet_memory_s2 = packet_memory_s2_grant_vector[1];

  //sgdma_rx/m_write saved-grant packet_memory/s2, which is an e_assign
  assign sgdma_rx_m_write_saved_grant_packet_memory_s2 = packet_memory_s2_arb_winner[1] && sgdma_rx_m_write_requests_packet_memory_s2;

  //packet_memory/s2 chosen-master double-vector, which is an e_assign
  assign packet_memory_s2_chosen_master_double_vector = {packet_memory_s2_master_qreq_vector, packet_memory_s2_master_qreq_vector} & ({~packet_memory_s2_master_qreq_vector, ~packet_memory_s2_master_qreq_vector} + packet_memory_s2_arb_addend);

  //stable onehot encoding of arb winner
  assign packet_memory_s2_arb_winner = (packet_memory_s2_allow_new_arb_cycle & | packet_memory_s2_grant_vector) ? packet_memory_s2_grant_vector : packet_memory_s2_saved_chosen_master_vector;

  //saved packet_memory_s2_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s2_saved_chosen_master_vector <= 0;
      else if (packet_memory_s2_allow_new_arb_cycle)
          packet_memory_s2_saved_chosen_master_vector <= |packet_memory_s2_grant_vector ? packet_memory_s2_grant_vector : packet_memory_s2_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign packet_memory_s2_grant_vector = {(packet_memory_s2_chosen_master_double_vector[1] | packet_memory_s2_chosen_master_double_vector[3]),
    (packet_memory_s2_chosen_master_double_vector[0] | packet_memory_s2_chosen_master_double_vector[2])};

  //packet_memory/s2 chosen master rotated left, which is an e_assign
  assign packet_memory_s2_chosen_master_rot_left = (packet_memory_s2_arb_winner << 1) ? (packet_memory_s2_arb_winner << 1) : 1;

  //packet_memory/s2's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s2_arb_addend <= 1;
      else if (|packet_memory_s2_grant_vector)
          packet_memory_s2_arb_addend <= packet_memory_s2_end_xfer? packet_memory_s2_chosen_master_rot_left : packet_memory_s2_grant_vector;
    end


  assign packet_memory_s2_chipselect = sgdma_rx_m_write_granted_packet_memory_s2 | sgdma_tx_m_read_granted_packet_memory_s2;
  //packet_memory_s2_firsttransfer first transaction, which is an e_assign
  assign packet_memory_s2_firsttransfer = packet_memory_s2_begins_xfer ? packet_memory_s2_unreg_firsttransfer : packet_memory_s2_reg_firsttransfer;

  //packet_memory_s2_unreg_firsttransfer first transaction, which is an e_assign
  assign packet_memory_s2_unreg_firsttransfer = ~(packet_memory_s2_slavearbiterlockenable & packet_memory_s2_any_continuerequest);

  //packet_memory_s2_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          packet_memory_s2_reg_firsttransfer <= 1'b1;
      else if (packet_memory_s2_begins_xfer)
          packet_memory_s2_reg_firsttransfer <= packet_memory_s2_unreg_firsttransfer;
    end


  //packet_memory_s2_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign packet_memory_s2_beginbursttransfer_internal = packet_memory_s2_begins_xfer;

  //packet_memory_s2_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign packet_memory_s2_arbitration_holdoff_internal = packet_memory_s2_begins_xfer & packet_memory_s2_firsttransfer;

  //packet_memory_s2_write assignment, which is an e_mux
  assign packet_memory_s2_write = sgdma_rx_m_write_granted_packet_memory_s2 & sgdma_rx_m_write_write;

  assign shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write = sgdma_rx_m_write_address_to_slave;
  //packet_memory_s2_address mux, which is an e_mux
  assign packet_memory_s2_address = (sgdma_rx_m_write_granted_packet_memory_s2)? (shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write >> 2) :
    (shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read >> 2);

  assign shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read = sgdma_tx_m_read_address_to_slave;
  //d1_packet_memory_s2_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_packet_memory_s2_end_xfer <= 1;
      else 
        d1_packet_memory_s2_end_xfer <= packet_memory_s2_end_xfer;
    end


  //packet_memory_s2_waits_for_read in a cycle, which is an e_mux
  assign packet_memory_s2_waits_for_read = packet_memory_s2_in_a_read_cycle & 0;

  //packet_memory_s2_in_a_read_cycle assignment, which is an e_assign
  assign packet_memory_s2_in_a_read_cycle = sgdma_tx_m_read_granted_packet_memory_s2 & sgdma_tx_m_read_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = packet_memory_s2_in_a_read_cycle;

  //packet_memory_s2_waits_for_write in a cycle, which is an e_mux
  assign packet_memory_s2_waits_for_write = packet_memory_s2_in_a_write_cycle & 0;

  //packet_memory_s2_in_a_write_cycle assignment, which is an e_assign
  assign packet_memory_s2_in_a_write_cycle = sgdma_rx_m_write_granted_packet_memory_s2 & sgdma_rx_m_write_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = packet_memory_s2_in_a_write_cycle;

  assign wait_for_packet_memory_s2_counter = 0;
  //packet_memory_s2_byteenable byte enable port mux, which is an e_mux
  assign packet_memory_s2_byteenable = (sgdma_rx_m_write_granted_packet_memory_s2)? sgdma_rx_m_write_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //packet_memory/s2 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_m_write_granted_packet_memory_s2 + sgdma_tx_m_read_granted_packet_memory_s2 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_m_write_saved_grant_packet_memory_s2 + sgdma_tx_m_read_saved_grant_packet_memory_s2 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_clock_crossing_ddr2_cpu_m1_to_pipeline_bridge_ddr2_s1_module (
                                                                                   // inputs:
                                                                                    clear_fifo,
                                                                                    clk,
                                                                                    data_in,
                                                                                    read,
                                                                                    reset_n,
                                                                                    sync_reset,
                                                                                    write,

                                                                                   // outputs:
                                                                                    data_out,
                                                                                    empty,
                                                                                    fifo_contains_ones_n,
                                                                                    full
                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_ddr2_s1_arbitrator (
                                            // inputs:
                                             clk,
                                             clock_crossing_ddr2_cpu_m1_address_to_slave,
                                             clock_crossing_ddr2_cpu_m1_byteenable,
                                             clock_crossing_ddr2_cpu_m1_latency_counter,
                                             clock_crossing_ddr2_cpu_m1_nativeaddress,
                                             clock_crossing_ddr2_cpu_m1_read,
                                             clock_crossing_ddr2_cpu_m1_write,
                                             clock_crossing_ddr2_cpu_m1_writedata,
                                             pipeline_bridge_ddr2_s1_endofpacket,
                                             pipeline_bridge_ddr2_s1_readdata,
                                             pipeline_bridge_ddr2_s1_readdatavalid,
                                             pipeline_bridge_ddr2_s1_waitrequest,
                                             reset_n,

                                            // outputs:
                                             clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1,
                                             clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1,
                                             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1,
                                             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register,
                                             clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1,
                                             d1_pipeline_bridge_ddr2_s1_end_xfer,
                                             pipeline_bridge_ddr2_s1_address,
                                             pipeline_bridge_ddr2_s1_arbiterlock,
                                             pipeline_bridge_ddr2_s1_arbiterlock2,
                                             pipeline_bridge_ddr2_s1_burstcount,
                                             pipeline_bridge_ddr2_s1_byteenable,
                                             pipeline_bridge_ddr2_s1_chipselect,
                                             pipeline_bridge_ddr2_s1_debugaccess,
                                             pipeline_bridge_ddr2_s1_endofpacket_from_sa,
                                             pipeline_bridge_ddr2_s1_nativeaddress,
                                             pipeline_bridge_ddr2_s1_read,
                                             pipeline_bridge_ddr2_s1_readdata_from_sa,
                                             pipeline_bridge_ddr2_s1_reset_n,
                                             pipeline_bridge_ddr2_s1_waitrequest_from_sa,
                                             pipeline_bridge_ddr2_s1_write,
                                             pipeline_bridge_ddr2_s1_writedata
                                          )
;

  output           clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1;
  output           clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1;
  output           clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1;
  output           clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register;
  output           clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;
  output           d1_pipeline_bridge_ddr2_s1_end_xfer;
  output  [ 27: 0] pipeline_bridge_ddr2_s1_address;
  output           pipeline_bridge_ddr2_s1_arbiterlock;
  output           pipeline_bridge_ddr2_s1_arbiterlock2;
  output           pipeline_bridge_ddr2_s1_burstcount;
  output  [  3: 0] pipeline_bridge_ddr2_s1_byteenable;
  output           pipeline_bridge_ddr2_s1_chipselect;
  output           pipeline_bridge_ddr2_s1_debugaccess;
  output           pipeline_bridge_ddr2_s1_endofpacket_from_sa;
  output  [ 27: 0] pipeline_bridge_ddr2_s1_nativeaddress;
  output           pipeline_bridge_ddr2_s1_read;
  output  [ 31: 0] pipeline_bridge_ddr2_s1_readdata_from_sa;
  output           pipeline_bridge_ddr2_s1_reset_n;
  output           pipeline_bridge_ddr2_s1_waitrequest_from_sa;
  output           pipeline_bridge_ddr2_s1_write;
  output  [ 31: 0] pipeline_bridge_ddr2_s1_writedata;
  input            clk;
  input   [ 29: 0] clock_crossing_ddr2_cpu_m1_address_to_slave;
  input   [  3: 0] clock_crossing_ddr2_cpu_m1_byteenable;
  input            clock_crossing_ddr2_cpu_m1_latency_counter;
  input   [ 27: 0] clock_crossing_ddr2_cpu_m1_nativeaddress;
  input            clock_crossing_ddr2_cpu_m1_read;
  input            clock_crossing_ddr2_cpu_m1_write;
  input   [ 31: 0] clock_crossing_ddr2_cpu_m1_writedata;
  input            pipeline_bridge_ddr2_s1_endofpacket;
  input   [ 31: 0] pipeline_bridge_ddr2_s1_readdata;
  input            pipeline_bridge_ddr2_s1_readdatavalid;
  input            pipeline_bridge_ddr2_s1_waitrequest;
  input            reset_n;

  wire             clock_crossing_ddr2_cpu_m1_arbiterlock;
  wire             clock_crossing_ddr2_cpu_m1_arbiterlock2;
  wire             clock_crossing_ddr2_cpu_m1_continuerequest;
  wire             clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_rdv_fifo_empty_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_rdv_fifo_output_from_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register;
  wire             clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_saved_grant_pipeline_bridge_ddr2_s1;
  reg              d1_pipeline_bridge_ddr2_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 27: 0] pipeline_bridge_ddr2_s1_address;
  wire             pipeline_bridge_ddr2_s1_allgrants;
  wire             pipeline_bridge_ddr2_s1_allow_new_arb_cycle;
  wire             pipeline_bridge_ddr2_s1_any_bursting_master_saved_grant;
  wire             pipeline_bridge_ddr2_s1_any_continuerequest;
  wire             pipeline_bridge_ddr2_s1_arb_counter_enable;
  reg              pipeline_bridge_ddr2_s1_arb_share_counter;
  wire             pipeline_bridge_ddr2_s1_arb_share_counter_next_value;
  wire             pipeline_bridge_ddr2_s1_arb_share_set_values;
  wire             pipeline_bridge_ddr2_s1_arbiterlock;
  wire             pipeline_bridge_ddr2_s1_arbiterlock2;
  wire             pipeline_bridge_ddr2_s1_arbitration_holdoff_internal;
  wire             pipeline_bridge_ddr2_s1_beginbursttransfer_internal;
  wire             pipeline_bridge_ddr2_s1_begins_xfer;
  wire             pipeline_bridge_ddr2_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_ddr2_s1_byteenable;
  wire             pipeline_bridge_ddr2_s1_chipselect;
  wire             pipeline_bridge_ddr2_s1_debugaccess;
  wire             pipeline_bridge_ddr2_s1_end_xfer;
  wire             pipeline_bridge_ddr2_s1_endofpacket_from_sa;
  wire             pipeline_bridge_ddr2_s1_firsttransfer;
  wire             pipeline_bridge_ddr2_s1_grant_vector;
  wire             pipeline_bridge_ddr2_s1_in_a_read_cycle;
  wire             pipeline_bridge_ddr2_s1_in_a_write_cycle;
  wire             pipeline_bridge_ddr2_s1_master_qreq_vector;
  wire             pipeline_bridge_ddr2_s1_move_on_to_next_transaction;
  wire    [ 27: 0] pipeline_bridge_ddr2_s1_nativeaddress;
  wire             pipeline_bridge_ddr2_s1_non_bursting_master_requests;
  wire             pipeline_bridge_ddr2_s1_read;
  wire    [ 31: 0] pipeline_bridge_ddr2_s1_readdata_from_sa;
  wire             pipeline_bridge_ddr2_s1_readdatavalid_from_sa;
  reg              pipeline_bridge_ddr2_s1_reg_firsttransfer;
  wire             pipeline_bridge_ddr2_s1_reset_n;
  reg              pipeline_bridge_ddr2_s1_slavearbiterlockenable;
  wire             pipeline_bridge_ddr2_s1_slavearbiterlockenable2;
  wire             pipeline_bridge_ddr2_s1_unreg_firsttransfer;
  wire             pipeline_bridge_ddr2_s1_waitrequest_from_sa;
  wire             pipeline_bridge_ddr2_s1_waits_for_read;
  wire             pipeline_bridge_ddr2_s1_waits_for_write;
  wire             pipeline_bridge_ddr2_s1_write;
  wire    [ 31: 0] pipeline_bridge_ddr2_s1_writedata;
  wire    [ 29: 0] shifted_address_to_pipeline_bridge_ddr2_s1_from_clock_crossing_ddr2_cpu_m1;
  wire             wait_for_pipeline_bridge_ddr2_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pipeline_bridge_ddr2_s1_end_xfer;
    end


  assign pipeline_bridge_ddr2_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1));
  //assign pipeline_bridge_ddr2_s1_readdata_from_sa = pipeline_bridge_ddr2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_ddr2_s1_readdata_from_sa = pipeline_bridge_ddr2_s1_readdata;

  assign clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1 = (1) & (clock_crossing_ddr2_cpu_m1_read | clock_crossing_ddr2_cpu_m1_write);
  //assign pipeline_bridge_ddr2_s1_waitrequest_from_sa = pipeline_bridge_ddr2_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_ddr2_s1_waitrequest_from_sa = pipeline_bridge_ddr2_s1_waitrequest;

  //assign pipeline_bridge_ddr2_s1_readdatavalid_from_sa = pipeline_bridge_ddr2_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_ddr2_s1_readdatavalid_from_sa = pipeline_bridge_ddr2_s1_readdatavalid;

  //pipeline_bridge_ddr2_s1_arb_share_counter set values, which is an e_mux
  assign pipeline_bridge_ddr2_s1_arb_share_set_values = 1;

  //pipeline_bridge_ddr2_s1_non_bursting_master_requests mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_non_bursting_master_requests = clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1 |
    clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;

  //pipeline_bridge_ddr2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_any_bursting_master_saved_grant = 0;

  //pipeline_bridge_ddr2_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pipeline_bridge_ddr2_s1_arb_share_counter_next_value = pipeline_bridge_ddr2_s1_firsttransfer ? (pipeline_bridge_ddr2_s1_arb_share_set_values - 1) : |pipeline_bridge_ddr2_s1_arb_share_counter ? (pipeline_bridge_ddr2_s1_arb_share_counter - 1) : 0;

  //pipeline_bridge_ddr2_s1_allgrants all slave grants, which is an e_mux
  assign pipeline_bridge_ddr2_s1_allgrants = (|pipeline_bridge_ddr2_s1_grant_vector) |
    (|pipeline_bridge_ddr2_s1_grant_vector);

  //pipeline_bridge_ddr2_s1_end_xfer assignment, which is an e_assign
  assign pipeline_bridge_ddr2_s1_end_xfer = ~(pipeline_bridge_ddr2_s1_waits_for_read | pipeline_bridge_ddr2_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1 = pipeline_bridge_ddr2_s1_end_xfer & (~pipeline_bridge_ddr2_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pipeline_bridge_ddr2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pipeline_bridge_ddr2_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1 & pipeline_bridge_ddr2_s1_allgrants) | (end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1 & ~pipeline_bridge_ddr2_s1_non_bursting_master_requests);

  //pipeline_bridge_ddr2_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_s1_arb_share_counter <= 0;
      else if (pipeline_bridge_ddr2_s1_arb_counter_enable)
          pipeline_bridge_ddr2_s1_arb_share_counter <= pipeline_bridge_ddr2_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge_ddr2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_s1_slavearbiterlockenable <= 0;
      else if ((|pipeline_bridge_ddr2_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1) | (end_xfer_arb_share_counter_term_pipeline_bridge_ddr2_s1 & ~pipeline_bridge_ddr2_s1_non_bursting_master_requests))
          pipeline_bridge_ddr2_s1_slavearbiterlockenable <= |pipeline_bridge_ddr2_s1_arb_share_counter_next_value;
    end


  //clock_crossing_ddr2_cpu/m1 pipeline_bridge_ddr2/s1 arbiterlock, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_arbiterlock = pipeline_bridge_ddr2_s1_slavearbiterlockenable & clock_crossing_ddr2_cpu_m1_continuerequest;

  //pipeline_bridge_ddr2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pipeline_bridge_ddr2_s1_slavearbiterlockenable2 = |pipeline_bridge_ddr2_s1_arb_share_counter_next_value;

  //clock_crossing_ddr2_cpu/m1 pipeline_bridge_ddr2/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_arbiterlock2 = pipeline_bridge_ddr2_s1_slavearbiterlockenable2 & clock_crossing_ddr2_cpu_m1_continuerequest;

  //pipeline_bridge_ddr2_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pipeline_bridge_ddr2_s1_any_continuerequest = 1;

  //clock_crossing_ddr2_cpu_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_continuerequest = 1;

  assign clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1 = clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1 & ~((clock_crossing_ddr2_cpu_m1_read & ((clock_crossing_ddr2_cpu_m1_latency_counter != 0) | (1 < clock_crossing_ddr2_cpu_m1_latency_counter))));
  //unique name for pipeline_bridge_ddr2_s1_move_on_to_next_transaction, which is an e_assign
  assign pipeline_bridge_ddr2_s1_move_on_to_next_transaction = pipeline_bridge_ddr2_s1_readdatavalid_from_sa;

  //rdv_fifo_for_clock_crossing_ddr2_cpu_m1_to_pipeline_bridge_ddr2_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_clock_crossing_ddr2_cpu_m1_to_pipeline_bridge_ddr2_s1_module rdv_fifo_for_clock_crossing_ddr2_cpu_m1_to_pipeline_bridge_ddr2_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1),
      .data_out             (clock_crossing_ddr2_cpu_m1_rdv_fifo_output_from_pipeline_bridge_ddr2_s1),
      .empty                (),
      .fifo_contains_ones_n (clock_crossing_ddr2_cpu_m1_rdv_fifo_empty_pipeline_bridge_ddr2_s1),
      .full                 (),
      .read                 (pipeline_bridge_ddr2_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_ddr2_s1_waits_for_read)
    );

  assign clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register = ~clock_crossing_ddr2_cpu_m1_rdv_fifo_empty_pipeline_bridge_ddr2_s1;
  //local readdatavalid clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1, which is an e_mux
  assign clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1 = pipeline_bridge_ddr2_s1_readdatavalid_from_sa;

  //pipeline_bridge_ddr2_s1_writedata mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_writedata = clock_crossing_ddr2_cpu_m1_writedata;

  //assign pipeline_bridge_ddr2_s1_endofpacket_from_sa = pipeline_bridge_ddr2_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_ddr2_s1_endofpacket_from_sa = pipeline_bridge_ddr2_s1_endofpacket;

  //master is always granted when requested
  assign clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1 = clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1;

  //clock_crossing_ddr2_cpu/m1 saved-grant pipeline_bridge_ddr2/s1, which is an e_assign
  assign clock_crossing_ddr2_cpu_m1_saved_grant_pipeline_bridge_ddr2_s1 = clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;

  //allow new arb cycle for pipeline_bridge_ddr2/s1, which is an e_assign
  assign pipeline_bridge_ddr2_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pipeline_bridge_ddr2_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pipeline_bridge_ddr2_s1_master_qreq_vector = 1;

  //pipeline_bridge_ddr2_s1_reset_n assignment, which is an e_assign
  assign pipeline_bridge_ddr2_s1_reset_n = reset_n;

  assign pipeline_bridge_ddr2_s1_chipselect = clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1;
  //pipeline_bridge_ddr2_s1_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_ddr2_s1_firsttransfer = pipeline_bridge_ddr2_s1_begins_xfer ? pipeline_bridge_ddr2_s1_unreg_firsttransfer : pipeline_bridge_ddr2_s1_reg_firsttransfer;

  //pipeline_bridge_ddr2_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_ddr2_s1_unreg_firsttransfer = ~(pipeline_bridge_ddr2_s1_slavearbiterlockenable & pipeline_bridge_ddr2_s1_any_continuerequest);

  //pipeline_bridge_ddr2_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_s1_reg_firsttransfer <= 1'b1;
      else if (pipeline_bridge_ddr2_s1_begins_xfer)
          pipeline_bridge_ddr2_s1_reg_firsttransfer <= pipeline_bridge_ddr2_s1_unreg_firsttransfer;
    end


  //pipeline_bridge_ddr2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pipeline_bridge_ddr2_s1_beginbursttransfer_internal = pipeline_bridge_ddr2_s1_begins_xfer;

  //pipeline_bridge_ddr2_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pipeline_bridge_ddr2_s1_arbitration_holdoff_internal = pipeline_bridge_ddr2_s1_begins_xfer & pipeline_bridge_ddr2_s1_firsttransfer;

  //pipeline_bridge_ddr2_s1_read assignment, which is an e_mux
  assign pipeline_bridge_ddr2_s1_read = clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1 & clock_crossing_ddr2_cpu_m1_read;

  //pipeline_bridge_ddr2_s1_write assignment, which is an e_mux
  assign pipeline_bridge_ddr2_s1_write = clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1 & clock_crossing_ddr2_cpu_m1_write;

  assign shifted_address_to_pipeline_bridge_ddr2_s1_from_clock_crossing_ddr2_cpu_m1 = clock_crossing_ddr2_cpu_m1_address_to_slave;
  //pipeline_bridge_ddr2_s1_address mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_address = shifted_address_to_pipeline_bridge_ddr2_s1_from_clock_crossing_ddr2_cpu_m1 >> 2;

  //slaveid pipeline_bridge_ddr2_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_nativeaddress = clock_crossing_ddr2_cpu_m1_nativeaddress;

  //d1_pipeline_bridge_ddr2_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pipeline_bridge_ddr2_s1_end_xfer <= 1;
      else 
        d1_pipeline_bridge_ddr2_s1_end_xfer <= pipeline_bridge_ddr2_s1_end_xfer;
    end


  //pipeline_bridge_ddr2_s1_waits_for_read in a cycle, which is an e_mux
  assign pipeline_bridge_ddr2_s1_waits_for_read = pipeline_bridge_ddr2_s1_in_a_read_cycle & pipeline_bridge_ddr2_s1_waitrequest_from_sa;

  //pipeline_bridge_ddr2_s1_in_a_read_cycle assignment, which is an e_assign
  assign pipeline_bridge_ddr2_s1_in_a_read_cycle = clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1 & clock_crossing_ddr2_cpu_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pipeline_bridge_ddr2_s1_in_a_read_cycle;

  //pipeline_bridge_ddr2_s1_waits_for_write in a cycle, which is an e_mux
  assign pipeline_bridge_ddr2_s1_waits_for_write = pipeline_bridge_ddr2_s1_in_a_write_cycle & pipeline_bridge_ddr2_s1_waitrequest_from_sa;

  //pipeline_bridge_ddr2_s1_in_a_write_cycle assignment, which is an e_assign
  assign pipeline_bridge_ddr2_s1_in_a_write_cycle = clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1 & clock_crossing_ddr2_cpu_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pipeline_bridge_ddr2_s1_in_a_write_cycle;

  assign wait_for_pipeline_bridge_ddr2_s1_counter = 0;
  //pipeline_bridge_ddr2_s1_byteenable byte enable port mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_byteenable = (clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1)? clock_crossing_ddr2_cpu_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_burstcount = 1;

  //pipeline_bridge_ddr2/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pipeline_bridge_ddr2_s1_arbiterlock = clock_crossing_ddr2_cpu_m1_arbiterlock;

  //pipeline_bridge_ddr2/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pipeline_bridge_ddr2_s1_arbiterlock2 = clock_crossing_ddr2_cpu_m1_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pipeline_bridge_ddr2_s1_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_ddr2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_module (
                                                                    // inputs:
                                                                     clear_fifo,
                                                                     clk,
                                                                     data_in,
                                                                     read,
                                                                     reset_n,
                                                                     sync_reset,
                                                                     write,

                                                                    // outputs:
                                                                     data_out,
                                                                     empty,
                                                                     fifo_contains_ones_n,
                                                                     full
                                                                  )
;

  output  [  2: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  2: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  2: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  2: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  2: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  2: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  2: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  2: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  2: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  2: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  2: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  2: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  2: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  2: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  2: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  2: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  2: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  2: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  2: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  2: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  2: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  2: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  2: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  2: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  2: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  2: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  2: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  2: 0] p31_stage_31;
  wire             p3_full_3;
  wire    [  2: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  2: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  2: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  2: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  2: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  2: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  2: 0] p9_stage_9;
  reg     [  2: 0] stage_0;
  reg     [  2: 0] stage_1;
  reg     [  2: 0] stage_10;
  reg     [  2: 0] stage_11;
  reg     [  2: 0] stage_12;
  reg     [  2: 0] stage_13;
  reg     [  2: 0] stage_14;
  reg     [  2: 0] stage_15;
  reg     [  2: 0] stage_16;
  reg     [  2: 0] stage_17;
  reg     [  2: 0] stage_18;
  reg     [  2: 0] stage_19;
  reg     [  2: 0] stage_2;
  reg     [  2: 0] stage_20;
  reg     [  2: 0] stage_21;
  reg     [  2: 0] stage_22;
  reg     [  2: 0] stage_23;
  reg     [  2: 0] stage_24;
  reg     [  2: 0] stage_25;
  reg     [  2: 0] stage_26;
  reg     [  2: 0] stage_27;
  reg     [  2: 0] stage_28;
  reg     [  2: 0] stage_29;
  reg     [  2: 0] stage_3;
  reg     [  2: 0] stage_30;
  reg     [  2: 0] stage_31;
  reg     [  2: 0] stage_4;
  reg     [  2: 0] stage_5;
  reg     [  2: 0] stage_6;
  reg     [  2: 0] stage_7;
  reg     [  2: 0] stage_8;
  reg     [  2: 0] stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_ddr2_m1_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_ddr2_s1_end_xfer,
                                             ddr2_s1_readdata_from_sa,
                                             ddr2_s1_waitrequest_n_from_sa,
                                             pipeline_bridge_ddr2_m1_address,
                                             pipeline_bridge_ddr2_m1_burstcount,
                                             pipeline_bridge_ddr2_m1_byteenable,
                                             pipeline_bridge_ddr2_m1_chipselect,
                                             pipeline_bridge_ddr2_m1_granted_ddr2_s1,
                                             pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1,
                                             pipeline_bridge_ddr2_m1_read,
                                             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1,
                                             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register,
                                             pipeline_bridge_ddr2_m1_requests_ddr2_s1,
                                             pipeline_bridge_ddr2_m1_write,
                                             pipeline_bridge_ddr2_m1_writedata,
                                             reset_n,

                                            // outputs:
                                             pipeline_bridge_ddr2_m1_address_to_slave,
                                             pipeline_bridge_ddr2_m1_latency_counter,
                                             pipeline_bridge_ddr2_m1_readdata,
                                             pipeline_bridge_ddr2_m1_readdatavalid,
                                             pipeline_bridge_ddr2_m1_waitrequest
                                          )
;

  output  [ 29: 0] pipeline_bridge_ddr2_m1_address_to_slave;
  output           pipeline_bridge_ddr2_m1_latency_counter;
  output  [ 31: 0] pipeline_bridge_ddr2_m1_readdata;
  output           pipeline_bridge_ddr2_m1_readdatavalid;
  output           pipeline_bridge_ddr2_m1_waitrequest;
  input            clk;
  input            d1_ddr2_s1_end_xfer;
  input   [255: 0] ddr2_s1_readdata_from_sa;
  input            ddr2_s1_waitrequest_n_from_sa;
  input   [ 29: 0] pipeline_bridge_ddr2_m1_address;
  input            pipeline_bridge_ddr2_m1_burstcount;
  input   [  3: 0] pipeline_bridge_ddr2_m1_byteenable;
  input            pipeline_bridge_ddr2_m1_chipselect;
  input            pipeline_bridge_ddr2_m1_granted_ddr2_s1;
  input            pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1;
  input            pipeline_bridge_ddr2_m1_read;
  input            pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;
  input            pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register;
  input            pipeline_bridge_ddr2_m1_requests_ddr2_s1;
  input            pipeline_bridge_ddr2_m1_write;
  input   [ 31: 0] pipeline_bridge_ddr2_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire    [ 31: 0] ddr2_s1_readdata_from_sa_part_selected_by_negative_dbs;
  wire             empty_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo;
  wire             full_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo;
  wire             latency_load_value;
  wire             p1_pipeline_bridge_ddr2_m1_latency_counter;
  reg     [ 29: 0] pipeline_bridge_ddr2_m1_address_last_time;
  wire    [ 29: 0] pipeline_bridge_ddr2_m1_address_to_slave;
  reg              pipeline_bridge_ddr2_m1_burstcount_last_time;
  reg     [  3: 0] pipeline_bridge_ddr2_m1_byteenable_last_time;
  reg              pipeline_bridge_ddr2_m1_chipselect_last_time;
  wire             pipeline_bridge_ddr2_m1_is_granted_some_slave;
  reg              pipeline_bridge_ddr2_m1_latency_counter;
  reg              pipeline_bridge_ddr2_m1_read_but_no_slave_selected;
  reg              pipeline_bridge_ddr2_m1_read_last_time;
  wire    [ 31: 0] pipeline_bridge_ddr2_m1_readdata;
  wire             pipeline_bridge_ddr2_m1_readdatavalid;
  wire             pipeline_bridge_ddr2_m1_run;
  wire             pipeline_bridge_ddr2_m1_waitrequest;
  reg              pipeline_bridge_ddr2_m1_write_last_time;
  reg     [ 31: 0] pipeline_bridge_ddr2_m1_writedata_last_time;
  wire             pre_flush_pipeline_bridge_ddr2_m1_readdatavalid;
  wire             r_0;
  wire             read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo;
  wire    [  2: 0] selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output;
  wire    [  2: 0] selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1;
  wire             write_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1 | ~pipeline_bridge_ddr2_m1_requests_ddr2_s1) & (pipeline_bridge_ddr2_m1_granted_ddr2_s1 | ~pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1) & ((~pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1 | ~pipeline_bridge_ddr2_m1_chipselect | (1 & ddr2_s1_waitrequest_n_from_sa & pipeline_bridge_ddr2_m1_chipselect))) & ((~pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1 | ~pipeline_bridge_ddr2_m1_chipselect | (1 & ddr2_s1_waitrequest_n_from_sa & pipeline_bridge_ddr2_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign pipeline_bridge_ddr2_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign pipeline_bridge_ddr2_m1_address_to_slave = pipeline_bridge_ddr2_m1_address[29 : 0];

  //pipeline_bridge_ddr2_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_read_but_no_slave_selected <= 0;
      else 
        pipeline_bridge_ddr2_m1_read_but_no_slave_selected <= (pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect) & pipeline_bridge_ddr2_m1_run & ~pipeline_bridge_ddr2_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pipeline_bridge_ddr2_m1_is_granted_some_slave = pipeline_bridge_ddr2_m1_granted_ddr2_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pipeline_bridge_ddr2_m1_readdatavalid = pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pipeline_bridge_ddr2_m1_readdatavalid = pipeline_bridge_ddr2_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_ddr2_m1_readdatavalid;

  //Negative Dynamic Bus-sizing mux.
  //this mux selects the correct eighth of the 
  //wide data coming from the slave ddr2/s1 
  assign ddr2_s1_readdata_from_sa_part_selected_by_negative_dbs = ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 0))? ddr2_s1_readdata_from_sa[31 : 0] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 1))? ddr2_s1_readdata_from_sa[63 : 32] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 2))? ddr2_s1_readdata_from_sa[95 : 64] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 3))? ddr2_s1_readdata_from_sa[127 : 96] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 4))? ddr2_s1_readdata_from_sa[159 : 128] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 5))? ddr2_s1_readdata_from_sa[191 : 160] :
    ((selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 == 6))? ddr2_s1_readdata_from_sa[223 : 192] :
    ddr2_s1_readdata_from_sa[255 : 224];

  //read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo fifo read, which is an e_mux
  assign read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo = pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;

  //write_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo fifo write, which is an e_mux
  assign write_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo = (pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect) & pipeline_bridge_ddr2_m1_run & pipeline_bridge_ddr2_m1_requests_ddr2_s1;

  assign selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output_ddr2_s1 = selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output;
  //selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_module selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_ddr2_m1_address_to_slave[4 : 2]),
      .data_out             (selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo_output),
      .empty                (empty_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo),
      .fifo_contains_ones_n (),
      .full                 (full_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo),
      .read                 (read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (write_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo)
    );

  //pipeline_bridge_ddr2/m1 readdata mux, which is an e_mux
  assign pipeline_bridge_ddr2_m1_readdata = ddr2_s1_readdata_from_sa_part_selected_by_negative_dbs;

  //actual waitrequest port, which is an e_assign
  assign pipeline_bridge_ddr2_m1_waitrequest = ~pipeline_bridge_ddr2_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_latency_counter <= 0;
      else 
        pipeline_bridge_ddr2_m1_latency_counter <= p1_pipeline_bridge_ddr2_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pipeline_bridge_ddr2_m1_latency_counter = ((pipeline_bridge_ddr2_m1_run & (pipeline_bridge_ddr2_m1_read & pipeline_bridge_ddr2_m1_chipselect)))? latency_load_value :
    (pipeline_bridge_ddr2_m1_latency_counter)? pipeline_bridge_ddr2_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_ddr2_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_address_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_address_last_time <= pipeline_bridge_ddr2_m1_address;
    end


  //pipeline_bridge_ddr2/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pipeline_bridge_ddr2_m1_waitrequest & pipeline_bridge_ddr2_m1_chipselect;
    end


  //pipeline_bridge_ddr2_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_address != pipeline_bridge_ddr2_m1_address_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_chipselect_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_chipselect_last_time <= pipeline_bridge_ddr2_m1_chipselect;
    end


  //pipeline_bridge_ddr2_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_chipselect != pipeline_bridge_ddr2_m1_chipselect_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_burstcount_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_burstcount_last_time <= pipeline_bridge_ddr2_m1_burstcount;
    end


  //pipeline_bridge_ddr2_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_burstcount != pipeline_bridge_ddr2_m1_burstcount_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_byteenable_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_byteenable_last_time <= pipeline_bridge_ddr2_m1_byteenable;
    end


  //pipeline_bridge_ddr2_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_byteenable != pipeline_bridge_ddr2_m1_byteenable_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_read_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_read_last_time <= pipeline_bridge_ddr2_m1_read;
    end


  //pipeline_bridge_ddr2_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_read != pipeline_bridge_ddr2_m1_read_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_write_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_write_last_time <= pipeline_bridge_ddr2_m1_write;
    end


  //pipeline_bridge_ddr2_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_write != pipeline_bridge_ddr2_m1_write_last_time))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_ddr2_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_ddr2_m1_writedata_last_time <= 0;
      else 
        pipeline_bridge_ddr2_m1_writedata_last_time <= pipeline_bridge_ddr2_m1_writedata;
    end


  //pipeline_bridge_ddr2_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_ddr2_m1_writedata != pipeline_bridge_ddr2_m1_writedata_last_time) & (pipeline_bridge_ddr2_m1_write & pipeline_bridge_ddr2_m1_chipselect))
        begin
          $write("%0d ns: pipeline_bridge_ddr2_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end


  //selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo read when empty, which is an e_process
  always @(posedge clk)
    begin
      if (empty_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo & read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo)
        begin
          $write("%0d ns: pipeline_bridge_ddr2/m1 negative rdv fifo selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo: read AND empty.\n", $time);
          $stop;
        end
    end


  //selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo write when full, which is an e_process
  always @(posedge clk)
    begin
      if (full_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo & write_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo & ~read_selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo)
        begin
          $write("%0d ns: pipeline_bridge_ddr2/m1 negative rdv fifo selecto_nrdv_pipeline_bridge_ddr2_m1_3_ddr2_s1_fifo: write AND full.\n", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_ddr2_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pll_s1_arbitrator (
                           // inputs:
                            SS_OCT_SOPC_clock_0_out_address_to_slave,
                            SS_OCT_SOPC_clock_0_out_nativeaddress,
                            SS_OCT_SOPC_clock_0_out_read,
                            SS_OCT_SOPC_clock_0_out_write,
                            SS_OCT_SOPC_clock_0_out_writedata,
                            clk,
                            pll_s1_readdata,
                            pll_s1_resetrequest,
                            reset_n,

                           // outputs:
                            SS_OCT_SOPC_clock_0_out_granted_pll_s1,
                            SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1,
                            SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1,
                            SS_OCT_SOPC_clock_0_out_requests_pll_s1,
                            d1_pll_s1_end_xfer,
                            pll_s1_address,
                            pll_s1_chipselect,
                            pll_s1_read,
                            pll_s1_readdata_from_sa,
                            pll_s1_reset_n,
                            pll_s1_resetrequest_from_sa,
                            pll_s1_write,
                            pll_s1_writedata
                         )
;

  output           SS_OCT_SOPC_clock_0_out_granted_pll_s1;
  output           SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1;
  output           SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1;
  output           SS_OCT_SOPC_clock_0_out_requests_pll_s1;
  output           d1_pll_s1_end_xfer;
  output  [  2: 0] pll_s1_address;
  output           pll_s1_chipselect;
  output           pll_s1_read;
  output  [ 15: 0] pll_s1_readdata_from_sa;
  output           pll_s1_reset_n;
  output           pll_s1_resetrequest_from_sa;
  output           pll_s1_write;
  output  [ 15: 0] pll_s1_writedata;
  input   [  3: 0] SS_OCT_SOPC_clock_0_out_address_to_slave;
  input   [  2: 0] SS_OCT_SOPC_clock_0_out_nativeaddress;
  input            SS_OCT_SOPC_clock_0_out_read;
  input            SS_OCT_SOPC_clock_0_out_write;
  input   [ 15: 0] SS_OCT_SOPC_clock_0_out_writedata;
  input            clk;
  input   [ 15: 0] pll_s1_readdata;
  input            pll_s1_resetrequest;
  input            reset_n;

  wire             SS_OCT_SOPC_clock_0_out_arbiterlock;
  wire             SS_OCT_SOPC_clock_0_out_arbiterlock2;
  wire             SS_OCT_SOPC_clock_0_out_continuerequest;
  wire             SS_OCT_SOPC_clock_0_out_granted_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_requests_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_saved_grant_pll_s1;
  reg              d1_pll_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pll_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_allgrants;
  wire             pll_s1_allow_new_arb_cycle;
  wire             pll_s1_any_bursting_master_saved_grant;
  wire             pll_s1_any_continuerequest;
  wire             pll_s1_arb_counter_enable;
  reg              pll_s1_arb_share_counter;
  wire             pll_s1_arb_share_counter_next_value;
  wire             pll_s1_arb_share_set_values;
  wire             pll_s1_beginbursttransfer_internal;
  wire             pll_s1_begins_xfer;
  wire             pll_s1_chipselect;
  wire             pll_s1_end_xfer;
  wire             pll_s1_firsttransfer;
  wire             pll_s1_grant_vector;
  wire             pll_s1_in_a_read_cycle;
  wire             pll_s1_in_a_write_cycle;
  wire             pll_s1_master_qreq_vector;
  wire             pll_s1_non_bursting_master_requests;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  reg              pll_s1_reg_firsttransfer;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest_from_sa;
  reg              pll_s1_slavearbiterlockenable;
  wire             pll_s1_slavearbiterlockenable2;
  wire             pll_s1_unreg_firsttransfer;
  wire             pll_s1_waits_for_read;
  wire             pll_s1_waits_for_write;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             wait_for_pll_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pll_s1_end_xfer;
    end


  assign pll_s1_begins_xfer = ~d1_reasons_to_wait & ((SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1));
  //assign pll_s1_readdata_from_sa = pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_readdata_from_sa = pll_s1_readdata;

  assign SS_OCT_SOPC_clock_0_out_requests_pll_s1 = (1) & (SS_OCT_SOPC_clock_0_out_read | SS_OCT_SOPC_clock_0_out_write);
  //pll_s1_arb_share_counter set values, which is an e_mux
  assign pll_s1_arb_share_set_values = 1;

  //pll_s1_non_bursting_master_requests mux, which is an e_mux
  assign pll_s1_non_bursting_master_requests = SS_OCT_SOPC_clock_0_out_requests_pll_s1;

  //pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pll_s1_any_bursting_master_saved_grant = 0;

  //pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pll_s1_arb_share_counter_next_value = pll_s1_firsttransfer ? (pll_s1_arb_share_set_values - 1) : |pll_s1_arb_share_counter ? (pll_s1_arb_share_counter - 1) : 0;

  //pll_s1_allgrants all slave grants, which is an e_mux
  assign pll_s1_allgrants = |pll_s1_grant_vector;

  //pll_s1_end_xfer assignment, which is an e_assign
  assign pll_s1_end_xfer = ~(pll_s1_waits_for_read | pll_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pll_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pll_s1 = pll_s1_end_xfer & (~pll_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pll_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pll_s1 & pll_s1_allgrants) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests);

  //pll_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_arb_share_counter <= 0;
      else if (pll_s1_arb_counter_enable)
          pll_s1_arb_share_counter <= pll_s1_arb_share_counter_next_value;
    end


  //pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_slavearbiterlockenable <= 0;
      else if ((|pll_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pll_s1) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests))
          pll_s1_slavearbiterlockenable <= |pll_s1_arb_share_counter_next_value;
    end


  //SS_OCT_SOPC_clock_0/out pll/s1 arbiterlock, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_arbiterlock = pll_s1_slavearbiterlockenable & SS_OCT_SOPC_clock_0_out_continuerequest;

  //pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pll_s1_slavearbiterlockenable2 = |pll_s1_arb_share_counter_next_value;

  //SS_OCT_SOPC_clock_0/out pll/s1 arbiterlock2, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_arbiterlock2 = pll_s1_slavearbiterlockenable2 & SS_OCT_SOPC_clock_0_out_continuerequest;

  //pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pll_s1_any_continuerequest = 1;

  //SS_OCT_SOPC_clock_0_out_continuerequest continued request, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_continuerequest = 1;

  assign SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1 = SS_OCT_SOPC_clock_0_out_requests_pll_s1;
  //pll_s1_writedata mux, which is an e_mux
  assign pll_s1_writedata = SS_OCT_SOPC_clock_0_out_writedata;

  //master is always granted when requested
  assign SS_OCT_SOPC_clock_0_out_granted_pll_s1 = SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1;

  //SS_OCT_SOPC_clock_0/out saved-grant pll/s1, which is an e_assign
  assign SS_OCT_SOPC_clock_0_out_saved_grant_pll_s1 = SS_OCT_SOPC_clock_0_out_requests_pll_s1;

  //allow new arb cycle for pll/s1, which is an e_assign
  assign pll_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pll_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pll_s1_master_qreq_vector = 1;

  //pll_s1_reset_n assignment, which is an e_assign
  assign pll_s1_reset_n = reset_n;

  //assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest;

  assign pll_s1_chipselect = SS_OCT_SOPC_clock_0_out_granted_pll_s1;
  //pll_s1_firsttransfer first transaction, which is an e_assign
  assign pll_s1_firsttransfer = pll_s1_begins_xfer ? pll_s1_unreg_firsttransfer : pll_s1_reg_firsttransfer;

  //pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pll_s1_unreg_firsttransfer = ~(pll_s1_slavearbiterlockenable & pll_s1_any_continuerequest);

  //pll_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_reg_firsttransfer <= 1'b1;
      else if (pll_s1_begins_xfer)
          pll_s1_reg_firsttransfer <= pll_s1_unreg_firsttransfer;
    end


  //pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pll_s1_beginbursttransfer_internal = pll_s1_begins_xfer;

  //pll_s1_read assignment, which is an e_mux
  assign pll_s1_read = SS_OCT_SOPC_clock_0_out_granted_pll_s1 & SS_OCT_SOPC_clock_0_out_read;

  //pll_s1_write assignment, which is an e_mux
  assign pll_s1_write = SS_OCT_SOPC_clock_0_out_granted_pll_s1 & SS_OCT_SOPC_clock_0_out_write;

  //pll_s1_address mux, which is an e_mux
  assign pll_s1_address = SS_OCT_SOPC_clock_0_out_nativeaddress;

  //d1_pll_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pll_s1_end_xfer <= 1;
      else 
        d1_pll_s1_end_xfer <= pll_s1_end_xfer;
    end


  //pll_s1_waits_for_read in a cycle, which is an e_mux
  assign pll_s1_waits_for_read = pll_s1_in_a_read_cycle & pll_s1_begins_xfer;

  //pll_s1_in_a_read_cycle assignment, which is an e_assign
  assign pll_s1_in_a_read_cycle = SS_OCT_SOPC_clock_0_out_granted_pll_s1 & SS_OCT_SOPC_clock_0_out_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pll_s1_in_a_read_cycle;

  //pll_s1_waits_for_write in a cycle, which is an e_mux
  assign pll_s1_waits_for_write = pll_s1_in_a_write_cycle & 0;

  //pll_s1_in_a_write_cycle assignment, which is an e_assign
  assign pll_s1_in_a_write_cycle = SS_OCT_SOPC_clock_0_out_granted_pll_s1 & SS_OCT_SOPC_clock_0_out_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pll_s1_in_a_write_cycle;

  assign wait_for_pll_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pll/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_latency_counter,
                                  cpu_data_master_read,
                                  cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,
                                  sgdma_rx_csr_irq,
                                  sgdma_rx_csr_readdata,

                                 // outputs:
                                  cpu_data_master_granted_sgdma_rx_csr,
                                  cpu_data_master_qualified_request_sgdma_rx_csr,
                                  cpu_data_master_read_data_valid_sgdma_rx_csr,
                                  cpu_data_master_requests_sgdma_rx_csr,
                                  d1_sgdma_rx_csr_end_xfer,
                                  sgdma_rx_csr_address,
                                  sgdma_rx_csr_chipselect,
                                  sgdma_rx_csr_irq_from_sa,
                                  sgdma_rx_csr_read,
                                  sgdma_rx_csr_readdata_from_sa,
                                  sgdma_rx_csr_reset_n,
                                  sgdma_rx_csr_write,
                                  sgdma_rx_csr_writedata
                               )
;

  output           cpu_data_master_granted_sgdma_rx_csr;
  output           cpu_data_master_qualified_request_sgdma_rx_csr;
  output           cpu_data_master_read_data_valid_sgdma_rx_csr;
  output           cpu_data_master_requests_sgdma_rx_csr;
  output           d1_sgdma_rx_csr_end_xfer;
  output  [  3: 0] sgdma_rx_csr_address;
  output           sgdma_rx_csr_chipselect;
  output           sgdma_rx_csr_irq_from_sa;
  output           sgdma_rx_csr_read;
  output  [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  output           sgdma_rx_csr_reset_n;
  output           sgdma_rx_csr_write;
  output  [ 31: 0] sgdma_rx_csr_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            sgdma_rx_csr_irq;
  input   [ 31: 0] sgdma_rx_csr_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sgdma_rx_csr;
  wire             cpu_data_master_qualified_request_sgdma_rx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_rx_csr;
  wire             cpu_data_master_requests_sgdma_rx_csr;
  wire             cpu_data_master_saved_grant_sgdma_rx_csr;
  reg              d1_reasons_to_wait;
  reg              d1_sgdma_rx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_rx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_allgrants;
  wire             sgdma_rx_csr_allow_new_arb_cycle;
  wire             sgdma_rx_csr_any_bursting_master_saved_grant;
  wire             sgdma_rx_csr_any_continuerequest;
  wire             sgdma_rx_csr_arb_counter_enable;
  reg     [  1: 0] sgdma_rx_csr_arb_share_counter;
  wire    [  1: 0] sgdma_rx_csr_arb_share_counter_next_value;
  wire    [  1: 0] sgdma_rx_csr_arb_share_set_values;
  wire             sgdma_rx_csr_beginbursttransfer_internal;
  wire             sgdma_rx_csr_begins_xfer;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_end_xfer;
  wire             sgdma_rx_csr_firsttransfer;
  wire             sgdma_rx_csr_grant_vector;
  wire             sgdma_rx_csr_in_a_read_cycle;
  wire             sgdma_rx_csr_in_a_write_cycle;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_master_qreq_vector;
  wire             sgdma_rx_csr_non_bursting_master_requests;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  reg              sgdma_rx_csr_reg_firsttransfer;
  wire             sgdma_rx_csr_reset_n;
  reg              sgdma_rx_csr_slavearbiterlockenable;
  wire             sgdma_rx_csr_slavearbiterlockenable2;
  wire             sgdma_rx_csr_unreg_firsttransfer;
  wire             sgdma_rx_csr_waits_for_read;
  wire             sgdma_rx_csr_waits_for_write;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 30: 0] shifted_address_to_sgdma_rx_csr_from_cpu_data_master;
  wire             wait_for_sgdma_rx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_rx_csr_end_xfer;
    end


  assign sgdma_rx_csr_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sgdma_rx_csr));
  //assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata;

  assign cpu_data_master_requests_sgdma_rx_csr = ({cpu_data_master_address_to_slave[30 : 6] , 6'b0} == 31'h481128c0) & (cpu_data_master_read | cpu_data_master_write);
  //sgdma_rx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_rx_csr_arb_share_set_values = 1;

  //sgdma_rx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_rx_csr_non_bursting_master_requests = cpu_data_master_requests_sgdma_rx_csr;

  //sgdma_rx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_rx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_rx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_rx_csr_arb_share_counter_next_value = sgdma_rx_csr_firsttransfer ? (sgdma_rx_csr_arb_share_set_values - 1) : |sgdma_rx_csr_arb_share_counter ? (sgdma_rx_csr_arb_share_counter - 1) : 0;

  //sgdma_rx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_rx_csr_allgrants = |sgdma_rx_csr_grant_vector;

  //sgdma_rx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_rx_csr_end_xfer = ~(sgdma_rx_csr_waits_for_read | sgdma_rx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_rx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_rx_csr = sgdma_rx_csr_end_xfer & (~sgdma_rx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_rx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_rx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_rx_csr & sgdma_rx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests);

  //sgdma_rx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_arb_share_counter <= 0;
      else if (sgdma_rx_csr_arb_counter_enable)
          sgdma_rx_csr_arb_share_counter <= sgdma_rx_csr_arb_share_counter_next_value;
    end


  //sgdma_rx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_rx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_rx_csr) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests))
          sgdma_rx_csr_slavearbiterlockenable <= |sgdma_rx_csr_arb_share_counter_next_value;
    end


  //cpu/data_master sgdma_rx/csr arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sgdma_rx_csr_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sgdma_rx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_rx_csr_slavearbiterlockenable2 = |sgdma_rx_csr_arb_share_counter_next_value;

  //cpu/data_master sgdma_rx/csr arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sgdma_rx_csr_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sgdma_rx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_rx_csr_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sgdma_rx_csr = cpu_data_master_requests_sgdma_rx_csr & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sgdma_rx_csr, which is an e_mux
  assign cpu_data_master_read_data_valid_sgdma_rx_csr = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read & ~sgdma_rx_csr_waits_for_read;

  //sgdma_rx_csr_writedata mux, which is an e_mux
  assign sgdma_rx_csr_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_sgdma_rx_csr = cpu_data_master_qualified_request_sgdma_rx_csr;

  //cpu/data_master saved-grant sgdma_rx/csr, which is an e_assign
  assign cpu_data_master_saved_grant_sgdma_rx_csr = cpu_data_master_requests_sgdma_rx_csr;

  //allow new arb cycle for sgdma_rx/csr, which is an e_assign
  assign sgdma_rx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_rx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_rx_csr_master_qreq_vector = 1;

  //sgdma_rx_csr_reset_n assignment, which is an e_assign
  assign sgdma_rx_csr_reset_n = reset_n;

  assign sgdma_rx_csr_chipselect = cpu_data_master_granted_sgdma_rx_csr;
  //sgdma_rx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_firsttransfer = sgdma_rx_csr_begins_xfer ? sgdma_rx_csr_unreg_firsttransfer : sgdma_rx_csr_reg_firsttransfer;

  //sgdma_rx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_unreg_firsttransfer = ~(sgdma_rx_csr_slavearbiterlockenable & sgdma_rx_csr_any_continuerequest);

  //sgdma_rx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_rx_csr_begins_xfer)
          sgdma_rx_csr_reg_firsttransfer <= sgdma_rx_csr_unreg_firsttransfer;
    end


  //sgdma_rx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_rx_csr_beginbursttransfer_internal = sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_read assignment, which is an e_mux
  assign sgdma_rx_csr_read = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read;

  //sgdma_rx_csr_write assignment, which is an e_mux
  assign sgdma_rx_csr_write = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_write;

  assign shifted_address_to_sgdma_rx_csr_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sgdma_rx_csr_address mux, which is an e_mux
  assign sgdma_rx_csr_address = shifted_address_to_sgdma_rx_csr_from_cpu_data_master >> 2;

  //d1_sgdma_rx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_rx_csr_end_xfer <= 1;
      else 
        d1_sgdma_rx_csr_end_xfer <= sgdma_rx_csr_end_xfer;
    end


  //sgdma_rx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_read = sgdma_rx_csr_in_a_read_cycle & sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_read_cycle = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_rx_csr_in_a_read_cycle;

  //sgdma_rx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_write = sgdma_rx_csr_in_a_write_cycle & 0;

  //sgdma_rx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_write_cycle = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_rx_csr_in_a_write_cycle;

  assign wait_for_sgdma_rx_csr_counter = 0;
  //assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_in_arbitrator (
                                // inputs:
                                 clk,
                                 reset_n,
                                 sgdma_rx_in_ready,
                                 tse_mac_receive_data,
                                 tse_mac_receive_empty,
                                 tse_mac_receive_endofpacket,
                                 tse_mac_receive_error,
                                 tse_mac_receive_startofpacket,
                                 tse_mac_receive_valid,

                                // outputs:
                                 sgdma_rx_in_data,
                                 sgdma_rx_in_empty,
                                 sgdma_rx_in_endofpacket,
                                 sgdma_rx_in_error,
                                 sgdma_rx_in_ready_from_sa,
                                 sgdma_rx_in_startofpacket,
                                 sgdma_rx_in_valid
                              )
;

  output  [ 31: 0] sgdma_rx_in_data;
  output  [  3: 0] sgdma_rx_in_empty;
  output           sgdma_rx_in_endofpacket;
  output  [  5: 0] sgdma_rx_in_error;
  output           sgdma_rx_in_ready_from_sa;
  output           sgdma_rx_in_startofpacket;
  output           sgdma_rx_in_valid;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  3: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  //mux sgdma_rx_in_data, which is an e_mux
  assign sgdma_rx_in_data = tse_mac_receive_data;

  //mux sgdma_rx_in_empty, which is an e_mux
  assign sgdma_rx_in_empty = tse_mac_receive_empty;

  //mux sgdma_rx_in_endofpacket, which is an e_mux
  assign sgdma_rx_in_endofpacket = tse_mac_receive_endofpacket;

  //mux sgdma_rx_in_error, which is an e_mux
  assign sgdma_rx_in_error = tse_mac_receive_error;

  //assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready;

  //mux sgdma_rx_in_startofpacket, which is an e_mux
  assign sgdma_rx_in_startofpacket = tse_mac_receive_startofpacket;

  //mux sgdma_rx_in_valid, which is an e_mux
  assign sgdma_rx_in_valid = tse_mac_receive_valid;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_descriptor_memory_s1_end_xfer,
                                              descriptor_memory_s1_readdata_from_sa,
                                              reset_n,
                                              sgdma_rx_descriptor_read_address,
                                              sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_read,
                                              sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_requests_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_rx_descriptor_read_address_to_slave,
                                              sgdma_rx_descriptor_read_latency_counter,
                                              sgdma_rx_descriptor_read_readdata,
                                              sgdma_rx_descriptor_read_readdatavalid,
                                              sgdma_rx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  output           sgdma_rx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_rx_descriptor_read_readdata;
  output           sgdma_rx_descriptor_read_readdatavalid;
  output           sgdma_rx_descriptor_read_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address;
  input            sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_read;
  input            sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_requests_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_rx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_rx_descriptor_read_readdatavalid;
  wire             r_0;
  reg     [ 31: 0] sgdma_rx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_is_granted_some_slave;
  reg              sgdma_rx_descriptor_read_latency_counter;
  reg              sgdma_rx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_rx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_run;
  wire             sgdma_rx_descriptor_read_waitrequest;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_requests_descriptor_memory_s1) & (sgdma_rx_descriptor_read_granted_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1) & ((~sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | ~(sgdma_rx_descriptor_read_read) | (1 & (sgdma_rx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_read_address_to_slave = {21'b10010000001000100011,
    sgdma_rx_descriptor_read_address[10 : 0]};

  //sgdma_rx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_rx_descriptor_read_read_but_no_slave_selected <= sgdma_rx_descriptor_read_read & sgdma_rx_descriptor_read_run & ~sgdma_rx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_rx_descriptor_read_is_granted_some_slave = sgdma_rx_descriptor_read_granted_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_rx_descriptor_read_readdatavalid;

  //sgdma_rx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_rx_descriptor_read_readdata = descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_read_waitrequest = ~sgdma_rx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_rx_descriptor_read_latency_counter <= p1_sgdma_rx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_rx_descriptor_read_latency_counter = ((sgdma_rx_descriptor_read_run & sgdma_rx_descriptor_read_read))? latency_load_value :
    (sgdma_rx_descriptor_read_latency_counter)? sgdma_rx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {sgdma_rx_descriptor_read_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_address_last_time <= sgdma_rx_descriptor_read_address;
    end


  //sgdma_rx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_read_waitrequest & (sgdma_rx_descriptor_read_read);
    end


  //sgdma_rx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_address != sgdma_rx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_read_last_time <= sgdma_rx_descriptor_read_read;
    end


  //sgdma_rx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_read != sgdma_rx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_descriptor_memory_s1_end_xfer,
                                               reset_n,
                                               sgdma_rx_descriptor_write_address,
                                               sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_write,
                                               sgdma_rx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_rx_descriptor_write_address_to_slave,
                                               sgdma_rx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  output           sgdma_rx_descriptor_write_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_write_address;
  input            sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_0;
  reg     [ 31: 0] sgdma_rx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_run;
  wire             sgdma_rx_descriptor_write_waitrequest;
  reg              sgdma_rx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_descriptor_write_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_requests_descriptor_memory_s1) & (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1) & ((~sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | ~(sgdma_rx_descriptor_write_write) | (1 & (sgdma_rx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_write_address_to_slave = {21'b10010000001000100011,
    sgdma_rx_descriptor_write_address[10 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_write_waitrequest = ~sgdma_rx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_address_last_time <= sgdma_rx_descriptor_write_address;
    end


  //sgdma_rx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_write_waitrequest & (sgdma_rx_descriptor_write_write);
    end


  //sgdma_rx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_address != sgdma_rx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_write_last_time <= sgdma_rx_descriptor_write_write;
    end


  //sgdma_rx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_write != sgdma_rx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_writedata_last_time <= sgdma_rx_descriptor_write_writedata;
    end


  //sgdma_rx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_writedata != sgdma_rx_descriptor_write_writedata_last_time) & sgdma_rx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_m_write_arbitrator (
                                     // inputs:
                                      clk,
                                      d1_onchip_memory_s1_end_xfer,
                                      d1_packet_memory_s2_end_xfer,
                                      reset_n,
                                      sgdma_rx_m_write_address,
                                      sgdma_rx_m_write_byteenable,
                                      sgdma_rx_m_write_granted_onchip_memory_s1,
                                      sgdma_rx_m_write_granted_packet_memory_s2,
                                      sgdma_rx_m_write_qualified_request_onchip_memory_s1,
                                      sgdma_rx_m_write_qualified_request_packet_memory_s2,
                                      sgdma_rx_m_write_requests_onchip_memory_s1,
                                      sgdma_rx_m_write_requests_packet_memory_s2,
                                      sgdma_rx_m_write_write,
                                      sgdma_rx_m_write_writedata,

                                     // outputs:
                                      sgdma_rx_m_write_address_to_slave,
                                      sgdma_rx_m_write_waitrequest
                                   )
;

  output  [ 31: 0] sgdma_rx_m_write_address_to_slave;
  output           sgdma_rx_m_write_waitrequest;
  input            clk;
  input            d1_onchip_memory_s1_end_xfer;
  input            d1_packet_memory_s2_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_granted_onchip_memory_s1;
  input            sgdma_rx_m_write_granted_packet_memory_s2;
  input            sgdma_rx_m_write_qualified_request_onchip_memory_s1;
  input            sgdma_rx_m_write_qualified_request_packet_memory_s2;
  input            sgdma_rx_m_write_requests_onchip_memory_s1;
  input            sgdma_rx_m_write_requests_packet_memory_s2;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_1;
  wire             r_2;
  reg     [ 31: 0] sgdma_rx_m_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  reg     [  3: 0] sgdma_rx_m_write_byteenable_last_time;
  wire             sgdma_rx_m_write_run;
  wire             sgdma_rx_m_write_waitrequest;
  reg              sgdma_rx_m_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_m_write_writedata_last_time;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_rx_m_write_qualified_request_onchip_memory_s1 | ~sgdma_rx_m_write_requests_onchip_memory_s1) & (sgdma_rx_m_write_granted_onchip_memory_s1 | ~sgdma_rx_m_write_qualified_request_onchip_memory_s1) & ((~sgdma_rx_m_write_qualified_request_onchip_memory_s1 | ~(sgdma_rx_m_write_write) | (1 & (sgdma_rx_m_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_m_write_run = r_1 & r_2;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (sgdma_rx_m_write_qualified_request_packet_memory_s2 | ~sgdma_rx_m_write_requests_packet_memory_s2) & (sgdma_rx_m_write_granted_packet_memory_s2 | ~sgdma_rx_m_write_qualified_request_packet_memory_s2) & ((~sgdma_rx_m_write_qualified_request_packet_memory_s2 | ~(sgdma_rx_m_write_write) | (1 & (sgdma_rx_m_write_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_m_write_address_to_slave = {11'b1001000000,
    sgdma_rx_m_write_address[20 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_m_write_waitrequest = ~sgdma_rx_m_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_m_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_address_last_time <= 0;
      else 
        sgdma_rx_m_write_address_last_time <= sgdma_rx_m_write_address;
    end


  //sgdma_rx/m_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_m_write_waitrequest & (sgdma_rx_m_write_write);
    end


  //sgdma_rx_m_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_address != sgdma_rx_m_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_byteenable_last_time <= 0;
      else 
        sgdma_rx_m_write_byteenable_last_time <= sgdma_rx_m_write_byteenable;
    end


  //sgdma_rx_m_write_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_byteenable != sgdma_rx_m_write_byteenable_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_write_last_time <= 0;
      else 
        sgdma_rx_m_write_write_last_time <= sgdma_rx_m_write_write;
    end


  //sgdma_rx_m_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_write != sgdma_rx_m_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_writedata_last_time <= 0;
      else 
        sgdma_rx_m_write_writedata_last_time <= sgdma_rx_m_write_writedata;
    end


  //sgdma_rx_m_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_writedata != sgdma_rx_m_write_writedata_last_time) & sgdma_rx_m_write_write)
        begin
          $write("%0d ns: sgdma_rx_m_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_latency_counter,
                                  cpu_data_master_read,
                                  cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,
                                  sgdma_tx_csr_irq,
                                  sgdma_tx_csr_readdata,

                                 // outputs:
                                  cpu_data_master_granted_sgdma_tx_csr,
                                  cpu_data_master_qualified_request_sgdma_tx_csr,
                                  cpu_data_master_read_data_valid_sgdma_tx_csr,
                                  cpu_data_master_requests_sgdma_tx_csr,
                                  d1_sgdma_tx_csr_end_xfer,
                                  sgdma_tx_csr_address,
                                  sgdma_tx_csr_chipselect,
                                  sgdma_tx_csr_irq_from_sa,
                                  sgdma_tx_csr_read,
                                  sgdma_tx_csr_readdata_from_sa,
                                  sgdma_tx_csr_reset_n,
                                  sgdma_tx_csr_write,
                                  sgdma_tx_csr_writedata
                               )
;

  output           cpu_data_master_granted_sgdma_tx_csr;
  output           cpu_data_master_qualified_request_sgdma_tx_csr;
  output           cpu_data_master_read_data_valid_sgdma_tx_csr;
  output           cpu_data_master_requests_sgdma_tx_csr;
  output           d1_sgdma_tx_csr_end_xfer;
  output  [  3: 0] sgdma_tx_csr_address;
  output           sgdma_tx_csr_chipselect;
  output           sgdma_tx_csr_irq_from_sa;
  output           sgdma_tx_csr_read;
  output  [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  output           sgdma_tx_csr_reset_n;
  output           sgdma_tx_csr_write;
  output  [ 31: 0] sgdma_tx_csr_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            sgdma_tx_csr_irq;
  input   [ 31: 0] sgdma_tx_csr_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sgdma_tx_csr;
  wire             cpu_data_master_qualified_request_sgdma_tx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_tx_csr;
  wire             cpu_data_master_requests_sgdma_tx_csr;
  wire             cpu_data_master_saved_grant_sgdma_tx_csr;
  reg              d1_reasons_to_wait;
  reg              d1_sgdma_tx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_tx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_allgrants;
  wire             sgdma_tx_csr_allow_new_arb_cycle;
  wire             sgdma_tx_csr_any_bursting_master_saved_grant;
  wire             sgdma_tx_csr_any_continuerequest;
  wire             sgdma_tx_csr_arb_counter_enable;
  reg     [  1: 0] sgdma_tx_csr_arb_share_counter;
  wire    [  1: 0] sgdma_tx_csr_arb_share_counter_next_value;
  wire    [  1: 0] sgdma_tx_csr_arb_share_set_values;
  wire             sgdma_tx_csr_beginbursttransfer_internal;
  wire             sgdma_tx_csr_begins_xfer;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_end_xfer;
  wire             sgdma_tx_csr_firsttransfer;
  wire             sgdma_tx_csr_grant_vector;
  wire             sgdma_tx_csr_in_a_read_cycle;
  wire             sgdma_tx_csr_in_a_write_cycle;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_master_qreq_vector;
  wire             sgdma_tx_csr_non_bursting_master_requests;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  reg              sgdma_tx_csr_reg_firsttransfer;
  wire             sgdma_tx_csr_reset_n;
  reg              sgdma_tx_csr_slavearbiterlockenable;
  wire             sgdma_tx_csr_slavearbiterlockenable2;
  wire             sgdma_tx_csr_unreg_firsttransfer;
  wire             sgdma_tx_csr_waits_for_read;
  wire             sgdma_tx_csr_waits_for_write;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 30: 0] shifted_address_to_sgdma_tx_csr_from_cpu_data_master;
  wire             wait_for_sgdma_tx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_tx_csr_end_xfer;
    end


  assign sgdma_tx_csr_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sgdma_tx_csr));
  //assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata;

  assign cpu_data_master_requests_sgdma_tx_csr = ({cpu_data_master_address_to_slave[30 : 6] , 6'b0} == 31'h48112880) & (cpu_data_master_read | cpu_data_master_write);
  //sgdma_tx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_tx_csr_arb_share_set_values = 1;

  //sgdma_tx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_tx_csr_non_bursting_master_requests = cpu_data_master_requests_sgdma_tx_csr;

  //sgdma_tx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_tx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_tx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_tx_csr_arb_share_counter_next_value = sgdma_tx_csr_firsttransfer ? (sgdma_tx_csr_arb_share_set_values - 1) : |sgdma_tx_csr_arb_share_counter ? (sgdma_tx_csr_arb_share_counter - 1) : 0;

  //sgdma_tx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_tx_csr_allgrants = |sgdma_tx_csr_grant_vector;

  //sgdma_tx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_tx_csr_end_xfer = ~(sgdma_tx_csr_waits_for_read | sgdma_tx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_tx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_tx_csr = sgdma_tx_csr_end_xfer & (~sgdma_tx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_tx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_tx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_tx_csr & sgdma_tx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests);

  //sgdma_tx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_arb_share_counter <= 0;
      else if (sgdma_tx_csr_arb_counter_enable)
          sgdma_tx_csr_arb_share_counter <= sgdma_tx_csr_arb_share_counter_next_value;
    end


  //sgdma_tx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_tx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_tx_csr) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests))
          sgdma_tx_csr_slavearbiterlockenable <= |sgdma_tx_csr_arb_share_counter_next_value;
    end


  //cpu/data_master sgdma_tx/csr arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sgdma_tx_csr_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sgdma_tx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_tx_csr_slavearbiterlockenable2 = |sgdma_tx_csr_arb_share_counter_next_value;

  //cpu/data_master sgdma_tx/csr arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sgdma_tx_csr_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sgdma_tx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_tx_csr_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sgdma_tx_csr = cpu_data_master_requests_sgdma_tx_csr & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sgdma_tx_csr, which is an e_mux
  assign cpu_data_master_read_data_valid_sgdma_tx_csr = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read & ~sgdma_tx_csr_waits_for_read;

  //sgdma_tx_csr_writedata mux, which is an e_mux
  assign sgdma_tx_csr_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_sgdma_tx_csr = cpu_data_master_qualified_request_sgdma_tx_csr;

  //cpu/data_master saved-grant sgdma_tx/csr, which is an e_assign
  assign cpu_data_master_saved_grant_sgdma_tx_csr = cpu_data_master_requests_sgdma_tx_csr;

  //allow new arb cycle for sgdma_tx/csr, which is an e_assign
  assign sgdma_tx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_tx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_tx_csr_master_qreq_vector = 1;

  //sgdma_tx_csr_reset_n assignment, which is an e_assign
  assign sgdma_tx_csr_reset_n = reset_n;

  assign sgdma_tx_csr_chipselect = cpu_data_master_granted_sgdma_tx_csr;
  //sgdma_tx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_firsttransfer = sgdma_tx_csr_begins_xfer ? sgdma_tx_csr_unreg_firsttransfer : sgdma_tx_csr_reg_firsttransfer;

  //sgdma_tx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_unreg_firsttransfer = ~(sgdma_tx_csr_slavearbiterlockenable & sgdma_tx_csr_any_continuerequest);

  //sgdma_tx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_tx_csr_begins_xfer)
          sgdma_tx_csr_reg_firsttransfer <= sgdma_tx_csr_unreg_firsttransfer;
    end


  //sgdma_tx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_tx_csr_beginbursttransfer_internal = sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_read assignment, which is an e_mux
  assign sgdma_tx_csr_read = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read;

  //sgdma_tx_csr_write assignment, which is an e_mux
  assign sgdma_tx_csr_write = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_write;

  assign shifted_address_to_sgdma_tx_csr_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sgdma_tx_csr_address mux, which is an e_mux
  assign sgdma_tx_csr_address = shifted_address_to_sgdma_tx_csr_from_cpu_data_master >> 2;

  //d1_sgdma_tx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_tx_csr_end_xfer <= 1;
      else 
        d1_sgdma_tx_csr_end_xfer <= sgdma_tx_csr_end_xfer;
    end


  //sgdma_tx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_read = sgdma_tx_csr_in_a_read_cycle & sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_read_cycle = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_tx_csr_in_a_read_cycle;

  //sgdma_tx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_write = sgdma_tx_csr_in_a_write_cycle & 0;

  //sgdma_tx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_write_cycle = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_tx_csr_in_a_write_cycle;

  assign wait_for_sgdma_tx_csr_counter = 0;
  //assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_descriptor_memory_s1_end_xfer,
                                              descriptor_memory_s1_readdata_from_sa,
                                              reset_n,
                                              sgdma_tx_descriptor_read_address,
                                              sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_read,
                                              sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_requests_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_tx_descriptor_read_address_to_slave,
                                              sgdma_tx_descriptor_read_latency_counter,
                                              sgdma_tx_descriptor_read_readdata,
                                              sgdma_tx_descriptor_read_readdatavalid,
                                              sgdma_tx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  output           sgdma_tx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_tx_descriptor_read_readdata;
  output           sgdma_tx_descriptor_read_readdatavalid;
  output           sgdma_tx_descriptor_read_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_read_address;
  input            sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_read;
  input            sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_requests_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_tx_descriptor_read_readdatavalid;
  wire             r_0;
  reg     [ 31: 0] sgdma_tx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_is_granted_some_slave;
  reg              sgdma_tx_descriptor_read_latency_counter;
  reg              sgdma_tx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_tx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_run;
  wire             sgdma_tx_descriptor_read_waitrequest;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_requests_descriptor_memory_s1) & (sgdma_tx_descriptor_read_granted_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1) & ((~sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | ~(sgdma_tx_descriptor_read_read) | (1 & (sgdma_tx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_read_address_to_slave = {21'b10010000001000100011,
    sgdma_tx_descriptor_read_address[10 : 0]};

  //sgdma_tx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_descriptor_read_read_but_no_slave_selected <= sgdma_tx_descriptor_read_read & sgdma_tx_descriptor_read_run & ~sgdma_tx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_descriptor_read_is_granted_some_slave = sgdma_tx_descriptor_read_granted_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_descriptor_read_readdatavalid;

  //sgdma_tx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_tx_descriptor_read_readdata = descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_read_waitrequest = ~sgdma_tx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_tx_descriptor_read_latency_counter <= p1_sgdma_tx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_descriptor_read_latency_counter = ((sgdma_tx_descriptor_read_run & sgdma_tx_descriptor_read_read))? latency_load_value :
    (sgdma_tx_descriptor_read_latency_counter)? sgdma_tx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {sgdma_tx_descriptor_read_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_address_last_time <= sgdma_tx_descriptor_read_address;
    end


  //sgdma_tx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_read_waitrequest & (sgdma_tx_descriptor_read_read);
    end


  //sgdma_tx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_address != sgdma_tx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_read_last_time <= sgdma_tx_descriptor_read_read;
    end


  //sgdma_tx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_read != sgdma_tx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_descriptor_memory_s1_end_xfer,
                                               reset_n,
                                               sgdma_tx_descriptor_write_address,
                                               sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_requests_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_write,
                                               sgdma_tx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_tx_descriptor_write_address_to_slave,
                                               sgdma_tx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  output           sgdma_tx_descriptor_write_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_write_address;
  input            sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_0;
  reg     [ 31: 0] sgdma_tx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_run;
  wire             sgdma_tx_descriptor_write_waitrequest;
  reg              sgdma_tx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_tx_descriptor_write_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_requests_descriptor_memory_s1) & (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1) & ((~sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 | ~(sgdma_tx_descriptor_write_write) | (1 & (sgdma_tx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_write_address_to_slave = {21'b10010000001000100011,
    sgdma_tx_descriptor_write_address[10 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_write_waitrequest = ~sgdma_tx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_address_last_time <= sgdma_tx_descriptor_write_address;
    end


  //sgdma_tx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_write_waitrequest & (sgdma_tx_descriptor_write_write);
    end


  //sgdma_tx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_address != sgdma_tx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_write_last_time <= sgdma_tx_descriptor_write_write;
    end


  //sgdma_tx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_write != sgdma_tx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_writedata_last_time <= sgdma_tx_descriptor_write_writedata;
    end


  //sgdma_tx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_writedata != sgdma_tx_descriptor_write_writedata_last_time) & sgdma_tx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_m_read_arbitrator (
                                    // inputs:
                                     clk,
                                     d1_onchip_memory_s1_end_xfer,
                                     d1_packet_memory_s2_end_xfer,
                                     onchip_memory_s1_readdata_from_sa,
                                     packet_memory_s2_readdata_from_sa,
                                     reset_n,
                                     sgdma_tx_m_read_address,
                                     sgdma_tx_m_read_granted_onchip_memory_s1,
                                     sgdma_tx_m_read_granted_packet_memory_s2,
                                     sgdma_tx_m_read_qualified_request_onchip_memory_s1,
                                     sgdma_tx_m_read_qualified_request_packet_memory_s2,
                                     sgdma_tx_m_read_read,
                                     sgdma_tx_m_read_read_data_valid_onchip_memory_s1,
                                     sgdma_tx_m_read_read_data_valid_packet_memory_s2,
                                     sgdma_tx_m_read_requests_onchip_memory_s1,
                                     sgdma_tx_m_read_requests_packet_memory_s2,

                                    // outputs:
                                     sgdma_tx_m_read_address_to_slave,
                                     sgdma_tx_m_read_latency_counter,
                                     sgdma_tx_m_read_readdata,
                                     sgdma_tx_m_read_readdatavalid,
                                     sgdma_tx_m_read_waitrequest
                                  )
;

  output  [ 31: 0] sgdma_tx_m_read_address_to_slave;
  output           sgdma_tx_m_read_latency_counter;
  output  [ 31: 0] sgdma_tx_m_read_readdata;
  output           sgdma_tx_m_read_readdatavalid;
  output           sgdma_tx_m_read_waitrequest;
  input            clk;
  input            d1_onchip_memory_s1_end_xfer;
  input            d1_packet_memory_s2_end_xfer;
  input   [ 31: 0] onchip_memory_s1_readdata_from_sa;
  input   [ 31: 0] packet_memory_s2_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_m_read_address;
  input            sgdma_tx_m_read_granted_onchip_memory_s1;
  input            sgdma_tx_m_read_granted_packet_memory_s2;
  input            sgdma_tx_m_read_qualified_request_onchip_memory_s1;
  input            sgdma_tx_m_read_qualified_request_packet_memory_s2;
  input            sgdma_tx_m_read_read;
  input            sgdma_tx_m_read_read_data_valid_onchip_memory_s1;
  input            sgdma_tx_m_read_read_data_valid_packet_memory_s2;
  input            sgdma_tx_m_read_requests_onchip_memory_s1;
  input            sgdma_tx_m_read_requests_packet_memory_s2;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_m_read_latency_counter;
  wire             pre_flush_sgdma_tx_m_read_readdatavalid;
  wire             r_1;
  wire             r_2;
  reg     [ 31: 0] sgdma_tx_m_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_is_granted_some_slave;
  reg              sgdma_tx_m_read_latency_counter;
  reg              sgdma_tx_m_read_read_but_no_slave_selected;
  reg              sgdma_tx_m_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_run;
  wire             sgdma_tx_m_read_waitrequest;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_tx_m_read_qualified_request_onchip_memory_s1 | ~sgdma_tx_m_read_requests_onchip_memory_s1) & (sgdma_tx_m_read_granted_onchip_memory_s1 | ~sgdma_tx_m_read_qualified_request_onchip_memory_s1) & ((~sgdma_tx_m_read_qualified_request_onchip_memory_s1 | ~(sgdma_tx_m_read_read) | (1 & (sgdma_tx_m_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_m_read_run = r_1 & r_2;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (sgdma_tx_m_read_qualified_request_packet_memory_s2 | ~sgdma_tx_m_read_requests_packet_memory_s2) & (sgdma_tx_m_read_granted_packet_memory_s2 | ~sgdma_tx_m_read_qualified_request_packet_memory_s2) & ((~sgdma_tx_m_read_qualified_request_packet_memory_s2 | ~(sgdma_tx_m_read_read) | (1 & (sgdma_tx_m_read_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_m_read_address_to_slave = {11'b1001000000,
    sgdma_tx_m_read_address[20 : 0]};

  //sgdma_tx_m_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_m_read_read_but_no_slave_selected <= sgdma_tx_m_read_read & sgdma_tx_m_read_run & ~sgdma_tx_m_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_m_read_is_granted_some_slave = sgdma_tx_m_read_granted_onchip_memory_s1 |
    sgdma_tx_m_read_granted_packet_memory_s2;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_data_valid_onchip_memory_s1 |
    sgdma_tx_m_read_read_data_valid_packet_memory_s2;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_m_read_readdatavalid |
    sgdma_tx_m_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_m_read_readdatavalid;

  //sgdma_tx/m_read readdata mux, which is an e_mux
  assign sgdma_tx_m_read_readdata = ({32 {~sgdma_tx_m_read_read_data_valid_onchip_memory_s1}} | onchip_memory_s1_readdata_from_sa) &
    ({32 {~sgdma_tx_m_read_read_data_valid_packet_memory_s2}} | packet_memory_s2_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_m_read_waitrequest = ~sgdma_tx_m_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_latency_counter <= 0;
      else 
        sgdma_tx_m_read_latency_counter <= p1_sgdma_tx_m_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_m_read_latency_counter = ((sgdma_tx_m_read_run & sgdma_tx_m_read_read))? latency_load_value :
    (sgdma_tx_m_read_latency_counter)? sgdma_tx_m_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {sgdma_tx_m_read_requests_onchip_memory_s1}} & 1) |
    ({1 {sgdma_tx_m_read_requests_packet_memory_s2}} & 1);


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_m_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_address_last_time <= 0;
      else 
        sgdma_tx_m_read_address_last_time <= sgdma_tx_m_read_address;
    end


  //sgdma_tx/m_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_m_read_waitrequest & (sgdma_tx_m_read_read);
    end


  //sgdma_tx_m_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_address != sgdma_tx_m_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_m_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_last_time <= 0;
      else 
        sgdma_tx_m_read_read_last_time <= sgdma_tx_m_read_read;
    end


  //sgdma_tx_m_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_read != sgdma_tx_m_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_out_arbitrator (
                                 // inputs:
                                  clk,
                                  reset_n,
                                  sgdma_tx_out_data,
                                  sgdma_tx_out_empty,
                                  sgdma_tx_out_endofpacket,
                                  sgdma_tx_out_error,
                                  sgdma_tx_out_startofpacket,
                                  sgdma_tx_out_valid,
                                  tse_mac_transmit_ready_from_sa,

                                 // outputs:
                                  sgdma_tx_out_ready
                               )
;

  output           sgdma_tx_out_ready;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready_from_sa;

  wire             sgdma_tx_out_ready;
  //mux sgdma_tx_out_ready, which is an e_mux
  assign sgdma_tx_out_ready = tse_mac_transmit_ready_from_sa;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sys_timer_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_latency_counter,
                                  cpu_data_master_read,
                                  cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,
                                  sys_timer_s1_irq,
                                  sys_timer_s1_readdata,

                                 // outputs:
                                  cpu_data_master_granted_sys_timer_s1,
                                  cpu_data_master_qualified_request_sys_timer_s1,
                                  cpu_data_master_read_data_valid_sys_timer_s1,
                                  cpu_data_master_requests_sys_timer_s1,
                                  d1_sys_timer_s1_end_xfer,
                                  sys_timer_s1_address,
                                  sys_timer_s1_chipselect,
                                  sys_timer_s1_irq_from_sa,
                                  sys_timer_s1_readdata_from_sa,
                                  sys_timer_s1_reset_n,
                                  sys_timer_s1_write_n,
                                  sys_timer_s1_writedata
                               )
;

  output           cpu_data_master_granted_sys_timer_s1;
  output           cpu_data_master_qualified_request_sys_timer_s1;
  output           cpu_data_master_read_data_valid_sys_timer_s1;
  output           cpu_data_master_requests_sys_timer_s1;
  output           d1_sys_timer_s1_end_xfer;
  output  [  2: 0] sys_timer_s1_address;
  output           sys_timer_s1_chipselect;
  output           sys_timer_s1_irq_from_sa;
  output  [ 15: 0] sys_timer_s1_readdata_from_sa;
  output           sys_timer_s1_reset_n;
  output           sys_timer_s1_write_n;
  output  [ 15: 0] sys_timer_s1_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            sys_timer_s1_irq;
  input   [ 15: 0] sys_timer_s1_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sys_timer_s1;
  wire             cpu_data_master_qualified_request_sys_timer_s1;
  wire             cpu_data_master_read_data_valid_sys_timer_s1;
  wire             cpu_data_master_requests_sys_timer_s1;
  wire             cpu_data_master_saved_grant_sys_timer_s1;
  reg              d1_reasons_to_wait;
  reg              d1_sys_timer_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sys_timer_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_sys_timer_s1_from_cpu_data_master;
  wire    [  2: 0] sys_timer_s1_address;
  wire             sys_timer_s1_allgrants;
  wire             sys_timer_s1_allow_new_arb_cycle;
  wire             sys_timer_s1_any_bursting_master_saved_grant;
  wire             sys_timer_s1_any_continuerequest;
  wire             sys_timer_s1_arb_counter_enable;
  reg     [  1: 0] sys_timer_s1_arb_share_counter;
  wire    [  1: 0] sys_timer_s1_arb_share_counter_next_value;
  wire    [  1: 0] sys_timer_s1_arb_share_set_values;
  wire             sys_timer_s1_beginbursttransfer_internal;
  wire             sys_timer_s1_begins_xfer;
  wire             sys_timer_s1_chipselect;
  wire             sys_timer_s1_end_xfer;
  wire             sys_timer_s1_firsttransfer;
  wire             sys_timer_s1_grant_vector;
  wire             sys_timer_s1_in_a_read_cycle;
  wire             sys_timer_s1_in_a_write_cycle;
  wire             sys_timer_s1_irq_from_sa;
  wire             sys_timer_s1_master_qreq_vector;
  wire             sys_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] sys_timer_s1_readdata_from_sa;
  reg              sys_timer_s1_reg_firsttransfer;
  wire             sys_timer_s1_reset_n;
  reg              sys_timer_s1_slavearbiterlockenable;
  wire             sys_timer_s1_slavearbiterlockenable2;
  wire             sys_timer_s1_unreg_firsttransfer;
  wire             sys_timer_s1_waits_for_read;
  wire             sys_timer_s1_waits_for_write;
  wire             sys_timer_s1_write_n;
  wire    [ 15: 0] sys_timer_s1_writedata;
  wire             wait_for_sys_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sys_timer_s1_end_xfer;
    end


  assign sys_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sys_timer_s1));
  //assign sys_timer_s1_readdata_from_sa = sys_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_timer_s1_readdata_from_sa = sys_timer_s1_readdata;

  assign cpu_data_master_requests_sys_timer_s1 = ({cpu_data_master_address_to_slave[30 : 5] , 5'b0} == 31'h48112600) & (cpu_data_master_read | cpu_data_master_write);
  //sys_timer_s1_arb_share_counter set values, which is an e_mux
  assign sys_timer_s1_arb_share_set_values = 1;

  //sys_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign sys_timer_s1_non_bursting_master_requests = cpu_data_master_requests_sys_timer_s1;

  //sys_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sys_timer_s1_any_bursting_master_saved_grant = 0;

  //sys_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sys_timer_s1_arb_share_counter_next_value = sys_timer_s1_firsttransfer ? (sys_timer_s1_arb_share_set_values - 1) : |sys_timer_s1_arb_share_counter ? (sys_timer_s1_arb_share_counter - 1) : 0;

  //sys_timer_s1_allgrants all slave grants, which is an e_mux
  assign sys_timer_s1_allgrants = |sys_timer_s1_grant_vector;

  //sys_timer_s1_end_xfer assignment, which is an e_assign
  assign sys_timer_s1_end_xfer = ~(sys_timer_s1_waits_for_read | sys_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sys_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sys_timer_s1 = sys_timer_s1_end_xfer & (~sys_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sys_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sys_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sys_timer_s1 & sys_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_sys_timer_s1 & ~sys_timer_s1_non_bursting_master_requests);

  //sys_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_timer_s1_arb_share_counter <= 0;
      else if (sys_timer_s1_arb_counter_enable)
          sys_timer_s1_arb_share_counter <= sys_timer_s1_arb_share_counter_next_value;
    end


  //sys_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_timer_s1_slavearbiterlockenable <= 0;
      else if ((|sys_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sys_timer_s1) | (end_xfer_arb_share_counter_term_sys_timer_s1 & ~sys_timer_s1_non_bursting_master_requests))
          sys_timer_s1_slavearbiterlockenable <= |sys_timer_s1_arb_share_counter_next_value;
    end


  //cpu/data_master sys_timer/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sys_timer_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sys_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sys_timer_s1_slavearbiterlockenable2 = |sys_timer_s1_arb_share_counter_next_value;

  //cpu/data_master sys_timer/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sys_timer_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sys_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sys_timer_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sys_timer_s1 = cpu_data_master_requests_sys_timer_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sys_timer_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_sys_timer_s1 = cpu_data_master_granted_sys_timer_s1 & cpu_data_master_read & ~sys_timer_s1_waits_for_read;

  //sys_timer_s1_writedata mux, which is an e_mux
  assign sys_timer_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_sys_timer_s1 = cpu_data_master_qualified_request_sys_timer_s1;

  //cpu/data_master saved-grant sys_timer/s1, which is an e_assign
  assign cpu_data_master_saved_grant_sys_timer_s1 = cpu_data_master_requests_sys_timer_s1;

  //allow new arb cycle for sys_timer/s1, which is an e_assign
  assign sys_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sys_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sys_timer_s1_master_qreq_vector = 1;

  //sys_timer_s1_reset_n assignment, which is an e_assign
  assign sys_timer_s1_reset_n = reset_n;

  assign sys_timer_s1_chipselect = cpu_data_master_granted_sys_timer_s1;
  //sys_timer_s1_firsttransfer first transaction, which is an e_assign
  assign sys_timer_s1_firsttransfer = sys_timer_s1_begins_xfer ? sys_timer_s1_unreg_firsttransfer : sys_timer_s1_reg_firsttransfer;

  //sys_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sys_timer_s1_unreg_firsttransfer = ~(sys_timer_s1_slavearbiterlockenable & sys_timer_s1_any_continuerequest);

  //sys_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_timer_s1_reg_firsttransfer <= 1'b1;
      else if (sys_timer_s1_begins_xfer)
          sys_timer_s1_reg_firsttransfer <= sys_timer_s1_unreg_firsttransfer;
    end


  //sys_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sys_timer_s1_beginbursttransfer_internal = sys_timer_s1_begins_xfer;

  //~sys_timer_s1_write_n assignment, which is an e_mux
  assign sys_timer_s1_write_n = ~(cpu_data_master_granted_sys_timer_s1 & cpu_data_master_write);

  assign shifted_address_to_sys_timer_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sys_timer_s1_address mux, which is an e_mux
  assign sys_timer_s1_address = shifted_address_to_sys_timer_s1_from_cpu_data_master >> 2;

  //d1_sys_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sys_timer_s1_end_xfer <= 1;
      else 
        d1_sys_timer_s1_end_xfer <= sys_timer_s1_end_xfer;
    end


  //sys_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign sys_timer_s1_waits_for_read = sys_timer_s1_in_a_read_cycle & sys_timer_s1_begins_xfer;

  //sys_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign sys_timer_s1_in_a_read_cycle = cpu_data_master_granted_sys_timer_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sys_timer_s1_in_a_read_cycle;

  //sys_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign sys_timer_s1_waits_for_write = sys_timer_s1_in_a_write_cycle & 0;

  //sys_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign sys_timer_s1_in_a_write_cycle = cpu_data_master_granted_sys_timer_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sys_timer_s1_in_a_write_cycle;

  assign wait_for_sys_timer_s1_counter = 0;
  //assign sys_timer_s1_irq_from_sa = sys_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_timer_s1_irq_from_sa = sys_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sys_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_data_master_address_to_slave,
                                         cpu_data_master_latency_counter,
                                         cpu_data_master_read,
                                         cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                         cpu_data_master_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         cpu_data_master_granted_sysid_control_slave,
                                         cpu_data_master_qualified_request_sysid_control_slave,
                                         cpu_data_master_read_data_valid_sysid_control_slave,
                                         cpu_data_master_requests_sysid_control_slave,
                                         d1_sysid_control_slave_end_xfer,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa
                                      )
;

  output           cpu_data_master_granted_sysid_control_slave;
  output           cpu_data_master_qualified_request_sysid_control_slave;
  output           cpu_data_master_read_data_valid_sysid_control_slave;
  output           cpu_data_master_requests_sysid_control_slave;
  output           d1_sysid_control_slave_end_xfer;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sysid_control_slave;
  wire             cpu_data_master_qualified_request_sysid_control_slave;
  wire             cpu_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_data_master_requests_sysid_control_slave;
  wire             cpu_data_master_saved_grant_sysid_control_slave;
  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_sysid_control_slave_from_cpu_data_master;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg     [  1: 0] sysid_control_slave_arb_share_counter;
  wire    [  1: 0] sysid_control_slave_arb_share_counter_next_value;
  wire    [  1: 0] sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign cpu_data_master_requests_sysid_control_slave = (({cpu_data_master_address_to_slave[30 : 3] , 3'b0} == 31'h48112800) & (cpu_data_master_read | cpu_data_master_write)) & cpu_data_master_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = cpu_data_master_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //cpu/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //cpu/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sysid_control_slave = cpu_data_master_requests_sysid_control_slave & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sysid_control_slave, which is an e_mux
  assign cpu_data_master_read_data_valid_sysid_control_slave = cpu_data_master_granted_sysid_control_slave & cpu_data_master_read & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign cpu_data_master_granted_sysid_control_slave = cpu_data_master_qualified_request_sysid_control_slave;

  //cpu/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_data_master_saved_grant_sysid_control_slave = cpu_data_master_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  assign shifted_address_to_sysid_control_slave_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = shifted_address_to_sysid_control_slave_from_cpu_data_master >> 2;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = cpu_data_master_granted_sysid_control_slave & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = cpu_data_master_granted_sysid_control_slave & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_control_port_arbitrator (
                                         // inputs:
                                          clk,
                                          cpu_data_master_address_to_slave,
                                          cpu_data_master_latency_counter,
                                          cpu_data_master_read,
                                          cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                          cpu_data_master_write,
                                          cpu_data_master_writedata,
                                          reset_n,
                                          tse_mac_control_port_readdata,
                                          tse_mac_control_port_waitrequest,

                                         // outputs:
                                          cpu_data_master_granted_tse_mac_control_port,
                                          cpu_data_master_qualified_request_tse_mac_control_port,
                                          cpu_data_master_read_data_valid_tse_mac_control_port,
                                          cpu_data_master_requests_tse_mac_control_port,
                                          d1_tse_mac_control_port_end_xfer,
                                          tse_mac_control_port_address,
                                          tse_mac_control_port_read,
                                          tse_mac_control_port_readdata_from_sa,
                                          tse_mac_control_port_reset,
                                          tse_mac_control_port_waitrequest_from_sa,
                                          tse_mac_control_port_write,
                                          tse_mac_control_port_writedata
                                       )
;

  output           cpu_data_master_granted_tse_mac_control_port;
  output           cpu_data_master_qualified_request_tse_mac_control_port;
  output           cpu_data_master_read_data_valid_tse_mac_control_port;
  output           cpu_data_master_requests_tse_mac_control_port;
  output           d1_tse_mac_control_port_end_xfer;
  output  [  7: 0] tse_mac_control_port_address;
  output           tse_mac_control_port_read;
  output  [ 31: 0] tse_mac_control_port_readdata_from_sa;
  output           tse_mac_control_port_reset;
  output           tse_mac_control_port_waitrequest_from_sa;
  output           tse_mac_control_port_write;
  output  [ 31: 0] tse_mac_control_port_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] tse_mac_control_port_readdata;
  input            tse_mac_control_port_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_tse_mac_control_port;
  wire             cpu_data_master_qualified_request_tse_mac_control_port;
  wire             cpu_data_master_read_data_valid_tse_mac_control_port;
  wire             cpu_data_master_requests_tse_mac_control_port;
  wire             cpu_data_master_saved_grant_tse_mac_control_port;
  reg              d1_reasons_to_wait;
  reg              d1_tse_mac_control_port_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tse_mac_control_port;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_tse_mac_control_port_from_cpu_data_master;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_allgrants;
  wire             tse_mac_control_port_allow_new_arb_cycle;
  wire             tse_mac_control_port_any_bursting_master_saved_grant;
  wire             tse_mac_control_port_any_continuerequest;
  wire             tse_mac_control_port_arb_counter_enable;
  reg     [  1: 0] tse_mac_control_port_arb_share_counter;
  wire    [  1: 0] tse_mac_control_port_arb_share_counter_next_value;
  wire    [  1: 0] tse_mac_control_port_arb_share_set_values;
  wire             tse_mac_control_port_beginbursttransfer_internal;
  wire             tse_mac_control_port_begins_xfer;
  wire             tse_mac_control_port_end_xfer;
  wire             tse_mac_control_port_firsttransfer;
  wire             tse_mac_control_port_grant_vector;
  wire             tse_mac_control_port_in_a_read_cycle;
  wire             tse_mac_control_port_in_a_write_cycle;
  wire             tse_mac_control_port_master_qreq_vector;
  wire             tse_mac_control_port_non_bursting_master_requests;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  reg              tse_mac_control_port_reg_firsttransfer;
  wire             tse_mac_control_port_reset;
  reg              tse_mac_control_port_slavearbiterlockenable;
  wire             tse_mac_control_port_slavearbiterlockenable2;
  wire             tse_mac_control_port_unreg_firsttransfer;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_waits_for_read;
  wire             tse_mac_control_port_waits_for_write;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire             wait_for_tse_mac_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tse_mac_control_port_end_xfer;
    end


  assign tse_mac_control_port_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_tse_mac_control_port));
  //assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata;

  assign cpu_data_master_requests_tse_mac_control_port = ({cpu_data_master_address_to_slave[30 : 10] , 10'b0} == 31'h48112000) & (cpu_data_master_read | cpu_data_master_write);
  //assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest;

  //tse_mac_control_port_arb_share_counter set values, which is an e_mux
  assign tse_mac_control_port_arb_share_set_values = 1;

  //tse_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  assign tse_mac_control_port_non_bursting_master_requests = cpu_data_master_requests_tse_mac_control_port;

  //tse_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign tse_mac_control_port_any_bursting_master_saved_grant = 0;

  //tse_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign tse_mac_control_port_arb_share_counter_next_value = tse_mac_control_port_firsttransfer ? (tse_mac_control_port_arb_share_set_values - 1) : |tse_mac_control_port_arb_share_counter ? (tse_mac_control_port_arb_share_counter - 1) : 0;

  //tse_mac_control_port_allgrants all slave grants, which is an e_mux
  assign tse_mac_control_port_allgrants = |tse_mac_control_port_grant_vector;

  //tse_mac_control_port_end_xfer assignment, which is an e_assign
  assign tse_mac_control_port_end_xfer = ~(tse_mac_control_port_waits_for_read | tse_mac_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_tse_mac_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tse_mac_control_port = tse_mac_control_port_end_xfer & (~tse_mac_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tse_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign tse_mac_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_tse_mac_control_port & tse_mac_control_port_allgrants) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests);

  //tse_mac_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_arb_share_counter <= 0;
      else if (tse_mac_control_port_arb_counter_enable)
          tse_mac_control_port_arb_share_counter <= tse_mac_control_port_arb_share_counter_next_value;
    end


  //tse_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_slavearbiterlockenable <= 0;
      else if ((|tse_mac_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_tse_mac_control_port) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests))
          tse_mac_control_port_slavearbiterlockenable <= |tse_mac_control_port_arb_share_counter_next_value;
    end


  //cpu/data_master tse_mac/control_port arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = tse_mac_control_port_slavearbiterlockenable & cpu_data_master_continuerequest;

  //tse_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tse_mac_control_port_slavearbiterlockenable2 = |tse_mac_control_port_arb_share_counter_next_value;

  //cpu/data_master tse_mac/control_port arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = tse_mac_control_port_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //tse_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tse_mac_control_port_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_tse_mac_control_port = cpu_data_master_requests_tse_mac_control_port & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_tse_mac_control_port, which is an e_mux
  assign cpu_data_master_read_data_valid_tse_mac_control_port = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read & ~tse_mac_control_port_waits_for_read;

  //tse_mac_control_port_writedata mux, which is an e_mux
  assign tse_mac_control_port_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_tse_mac_control_port = cpu_data_master_qualified_request_tse_mac_control_port;

  //cpu/data_master saved-grant tse_mac/control_port, which is an e_assign
  assign cpu_data_master_saved_grant_tse_mac_control_port = cpu_data_master_requests_tse_mac_control_port;

  //allow new arb cycle for tse_mac/control_port, which is an e_assign
  assign tse_mac_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tse_mac_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tse_mac_control_port_master_qreq_vector = 1;

  //~tse_mac_control_port_reset assignment, which is an e_assign
  assign tse_mac_control_port_reset = ~reset_n;

  //tse_mac_control_port_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_firsttransfer = tse_mac_control_port_begins_xfer ? tse_mac_control_port_unreg_firsttransfer : tse_mac_control_port_reg_firsttransfer;

  //tse_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_unreg_firsttransfer = ~(tse_mac_control_port_slavearbiterlockenable & tse_mac_control_port_any_continuerequest);

  //tse_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_reg_firsttransfer <= 1'b1;
      else if (tse_mac_control_port_begins_xfer)
          tse_mac_control_port_reg_firsttransfer <= tse_mac_control_port_unreg_firsttransfer;
    end


  //tse_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tse_mac_control_port_beginbursttransfer_internal = tse_mac_control_port_begins_xfer;

  //tse_mac_control_port_read assignment, which is an e_mux
  assign tse_mac_control_port_read = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read;

  //tse_mac_control_port_write assignment, which is an e_mux
  assign tse_mac_control_port_write = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_write;

  assign shifted_address_to_tse_mac_control_port_from_cpu_data_master = cpu_data_master_address_to_slave;
  //tse_mac_control_port_address mux, which is an e_mux
  assign tse_mac_control_port_address = shifted_address_to_tse_mac_control_port_from_cpu_data_master >> 2;

  //d1_tse_mac_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tse_mac_control_port_end_xfer <= 1;
      else 
        d1_tse_mac_control_port_end_xfer <= tse_mac_control_port_end_xfer;
    end


  //tse_mac_control_port_waits_for_read in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_read = tse_mac_control_port_in_a_read_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_read_cycle = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tse_mac_control_port_in_a_read_cycle;

  //tse_mac_control_port_waits_for_write in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_write = tse_mac_control_port_in_a_write_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_write_cycle = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tse_mac_control_port_in_a_write_cycle;

  assign wait_for_tse_mac_control_port_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tse_mac/control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_transmit_arbitrator (
                                     // inputs:
                                      clk,
                                      reset_n,
                                      sgdma_tx_out_data,
                                      sgdma_tx_out_empty,
                                      sgdma_tx_out_endofpacket,
                                      sgdma_tx_out_error,
                                      sgdma_tx_out_startofpacket,
                                      sgdma_tx_out_valid,
                                      tse_mac_transmit_ready,

                                     // outputs:
                                      tse_mac_transmit_data,
                                      tse_mac_transmit_empty,
                                      tse_mac_transmit_endofpacket,
                                      tse_mac_transmit_error,
                                      tse_mac_transmit_ready_from_sa,
                                      tse_mac_transmit_startofpacket,
                                      tse_mac_transmit_valid
                                   )
;

  output  [ 31: 0] tse_mac_transmit_data;
  output  [  1: 0] tse_mac_transmit_empty;
  output           tse_mac_transmit_endofpacket;
  output           tse_mac_transmit_error;
  output           tse_mac_transmit_ready_from_sa;
  output           tse_mac_transmit_startofpacket;
  output           tse_mac_transmit_valid;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready;

  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  //mux tse_mac_transmit_data, which is an e_mux
  assign tse_mac_transmit_data = sgdma_tx_out_data;

  //mux tse_mac_transmit_endofpacket, which is an e_mux
  assign tse_mac_transmit_endofpacket = sgdma_tx_out_endofpacket;

  //mux tse_mac_transmit_error, which is an e_mux
  assign tse_mac_transmit_error = sgdma_tx_out_error;

  //mux tse_mac_transmit_empty, which is an e_mux
  assign tse_mac_transmit_empty = sgdma_tx_out_empty;

  //assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready;

  //mux tse_mac_transmit_startofpacket, which is an e_mux
  assign tse_mac_transmit_startofpacket = sgdma_tx_out_startofpacket;

  //mux tse_mac_transmit_valid, which is an e_mux
  assign tse_mac_transmit_valid = sgdma_tx_out_valid;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_receive_arbitrator (
                                    // inputs:
                                     clk,
                                     reset_n,
                                     sgdma_rx_in_ready_from_sa,
                                     tse_mac_receive_data,
                                     tse_mac_receive_empty,
                                     tse_mac_receive_endofpacket,
                                     tse_mac_receive_error,
                                     tse_mac_receive_startofpacket,
                                     tse_mac_receive_valid,

                                    // outputs:
                                     tse_mac_receive_ready
                                  )
;

  output           tse_mac_receive_ready;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready_from_sa;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire             tse_mac_receive_ready;
  //mux tse_mac_receive_ready, which is an e_mux
  assign tse_mac_receive_ready = sgdma_rx_in_ready_from_sa;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module vol_recording_done_pio_s1_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                               cpu_data_master_write,
                                               reset_n,
                                               vol_recording_done_pio_s1_readdata,

                                              // outputs:
                                               cpu_data_master_granted_vol_recording_done_pio_s1,
                                               cpu_data_master_qualified_request_vol_recording_done_pio_s1,
                                               cpu_data_master_read_data_valid_vol_recording_done_pio_s1,
                                               cpu_data_master_requests_vol_recording_done_pio_s1,
                                               d1_vol_recording_done_pio_s1_end_xfer,
                                               vol_recording_done_pio_s1_address,
                                               vol_recording_done_pio_s1_readdata_from_sa,
                                               vol_recording_done_pio_s1_reset_n
                                            )
;

  output           cpu_data_master_granted_vol_recording_done_pio_s1;
  output           cpu_data_master_qualified_request_vol_recording_done_pio_s1;
  output           cpu_data_master_read_data_valid_vol_recording_done_pio_s1;
  output           cpu_data_master_requests_vol_recording_done_pio_s1;
  output           d1_vol_recording_done_pio_s1_end_xfer;
  output  [  1: 0] vol_recording_done_pio_s1_address;
  output           vol_recording_done_pio_s1_readdata_from_sa;
  output           vol_recording_done_pio_s1_reset_n;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input            reset_n;
  input            vol_recording_done_pio_s1_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_vol_recording_done_pio_s1;
  wire             cpu_data_master_qualified_request_vol_recording_done_pio_s1;
  wire             cpu_data_master_read_data_valid_vol_recording_done_pio_s1;
  wire             cpu_data_master_requests_vol_recording_done_pio_s1;
  wire             cpu_data_master_saved_grant_vol_recording_done_pio_s1;
  reg              d1_reasons_to_wait;
  reg              d1_vol_recording_done_pio_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_vol_recording_done_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_vol_recording_done_pio_s1_from_cpu_data_master;
  wire    [  1: 0] vol_recording_done_pio_s1_address;
  wire             vol_recording_done_pio_s1_allgrants;
  wire             vol_recording_done_pio_s1_allow_new_arb_cycle;
  wire             vol_recording_done_pio_s1_any_bursting_master_saved_grant;
  wire             vol_recording_done_pio_s1_any_continuerequest;
  wire             vol_recording_done_pio_s1_arb_counter_enable;
  reg     [  1: 0] vol_recording_done_pio_s1_arb_share_counter;
  wire    [  1: 0] vol_recording_done_pio_s1_arb_share_counter_next_value;
  wire    [  1: 0] vol_recording_done_pio_s1_arb_share_set_values;
  wire             vol_recording_done_pio_s1_beginbursttransfer_internal;
  wire             vol_recording_done_pio_s1_begins_xfer;
  wire             vol_recording_done_pio_s1_end_xfer;
  wire             vol_recording_done_pio_s1_firsttransfer;
  wire             vol_recording_done_pio_s1_grant_vector;
  wire             vol_recording_done_pio_s1_in_a_read_cycle;
  wire             vol_recording_done_pio_s1_in_a_write_cycle;
  wire             vol_recording_done_pio_s1_master_qreq_vector;
  wire             vol_recording_done_pio_s1_non_bursting_master_requests;
  wire             vol_recording_done_pio_s1_readdata_from_sa;
  reg              vol_recording_done_pio_s1_reg_firsttransfer;
  wire             vol_recording_done_pio_s1_reset_n;
  reg              vol_recording_done_pio_s1_slavearbiterlockenable;
  wire             vol_recording_done_pio_s1_slavearbiterlockenable2;
  wire             vol_recording_done_pio_s1_unreg_firsttransfer;
  wire             vol_recording_done_pio_s1_waits_for_read;
  wire             vol_recording_done_pio_s1_waits_for_write;
  wire             wait_for_vol_recording_done_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~vol_recording_done_pio_s1_end_xfer;
    end


  assign vol_recording_done_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_vol_recording_done_pio_s1));
  //assign vol_recording_done_pio_s1_readdata_from_sa = vol_recording_done_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign vol_recording_done_pio_s1_readdata_from_sa = vol_recording_done_pio_s1_readdata;

  assign cpu_data_master_requests_vol_recording_done_pio_s1 = (({cpu_data_master_address_to_slave[30 : 4] , 4'b0} == 31'h48112780) & (cpu_data_master_read | cpu_data_master_write)) & cpu_data_master_read;
  //vol_recording_done_pio_s1_arb_share_counter set values, which is an e_mux
  assign vol_recording_done_pio_s1_arb_share_set_values = 1;

  //vol_recording_done_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign vol_recording_done_pio_s1_non_bursting_master_requests = cpu_data_master_requests_vol_recording_done_pio_s1;

  //vol_recording_done_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign vol_recording_done_pio_s1_any_bursting_master_saved_grant = 0;

  //vol_recording_done_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign vol_recording_done_pio_s1_arb_share_counter_next_value = vol_recording_done_pio_s1_firsttransfer ? (vol_recording_done_pio_s1_arb_share_set_values - 1) : |vol_recording_done_pio_s1_arb_share_counter ? (vol_recording_done_pio_s1_arb_share_counter - 1) : 0;

  //vol_recording_done_pio_s1_allgrants all slave grants, which is an e_mux
  assign vol_recording_done_pio_s1_allgrants = |vol_recording_done_pio_s1_grant_vector;

  //vol_recording_done_pio_s1_end_xfer assignment, which is an e_assign
  assign vol_recording_done_pio_s1_end_xfer = ~(vol_recording_done_pio_s1_waits_for_read | vol_recording_done_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_vol_recording_done_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_vol_recording_done_pio_s1 = vol_recording_done_pio_s1_end_xfer & (~vol_recording_done_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //vol_recording_done_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign vol_recording_done_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_vol_recording_done_pio_s1 & vol_recording_done_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_vol_recording_done_pio_s1 & ~vol_recording_done_pio_s1_non_bursting_master_requests);

  //vol_recording_done_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_recording_done_pio_s1_arb_share_counter <= 0;
      else if (vol_recording_done_pio_s1_arb_counter_enable)
          vol_recording_done_pio_s1_arb_share_counter <= vol_recording_done_pio_s1_arb_share_counter_next_value;
    end


  //vol_recording_done_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_recording_done_pio_s1_slavearbiterlockenable <= 0;
      else if ((|vol_recording_done_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_vol_recording_done_pio_s1) | (end_xfer_arb_share_counter_term_vol_recording_done_pio_s1 & ~vol_recording_done_pio_s1_non_bursting_master_requests))
          vol_recording_done_pio_s1_slavearbiterlockenable <= |vol_recording_done_pio_s1_arb_share_counter_next_value;
    end


  //cpu/data_master vol_recording_done_pio/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = vol_recording_done_pio_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //vol_recording_done_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign vol_recording_done_pio_s1_slavearbiterlockenable2 = |vol_recording_done_pio_s1_arb_share_counter_next_value;

  //cpu/data_master vol_recording_done_pio/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = vol_recording_done_pio_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //vol_recording_done_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign vol_recording_done_pio_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_vol_recording_done_pio_s1 = cpu_data_master_requests_vol_recording_done_pio_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_vol_recording_done_pio_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_vol_recording_done_pio_s1 = cpu_data_master_granted_vol_recording_done_pio_s1 & cpu_data_master_read & ~vol_recording_done_pio_s1_waits_for_read;

  //master is always granted when requested
  assign cpu_data_master_granted_vol_recording_done_pio_s1 = cpu_data_master_qualified_request_vol_recording_done_pio_s1;

  //cpu/data_master saved-grant vol_recording_done_pio/s1, which is an e_assign
  assign cpu_data_master_saved_grant_vol_recording_done_pio_s1 = cpu_data_master_requests_vol_recording_done_pio_s1;

  //allow new arb cycle for vol_recording_done_pio/s1, which is an e_assign
  assign vol_recording_done_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign vol_recording_done_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign vol_recording_done_pio_s1_master_qreq_vector = 1;

  //vol_recording_done_pio_s1_reset_n assignment, which is an e_assign
  assign vol_recording_done_pio_s1_reset_n = reset_n;

  //vol_recording_done_pio_s1_firsttransfer first transaction, which is an e_assign
  assign vol_recording_done_pio_s1_firsttransfer = vol_recording_done_pio_s1_begins_xfer ? vol_recording_done_pio_s1_unreg_firsttransfer : vol_recording_done_pio_s1_reg_firsttransfer;

  //vol_recording_done_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign vol_recording_done_pio_s1_unreg_firsttransfer = ~(vol_recording_done_pio_s1_slavearbiterlockenable & vol_recording_done_pio_s1_any_continuerequest);

  //vol_recording_done_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_recording_done_pio_s1_reg_firsttransfer <= 1'b1;
      else if (vol_recording_done_pio_s1_begins_xfer)
          vol_recording_done_pio_s1_reg_firsttransfer <= vol_recording_done_pio_s1_unreg_firsttransfer;
    end


  //vol_recording_done_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign vol_recording_done_pio_s1_beginbursttransfer_internal = vol_recording_done_pio_s1_begins_xfer;

  assign shifted_address_to_vol_recording_done_pio_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //vol_recording_done_pio_s1_address mux, which is an e_mux
  assign vol_recording_done_pio_s1_address = shifted_address_to_vol_recording_done_pio_s1_from_cpu_data_master >> 2;

  //d1_vol_recording_done_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_vol_recording_done_pio_s1_end_xfer <= 1;
      else 
        d1_vol_recording_done_pio_s1_end_xfer <= vol_recording_done_pio_s1_end_xfer;
    end


  //vol_recording_done_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign vol_recording_done_pio_s1_waits_for_read = vol_recording_done_pio_s1_in_a_read_cycle & vol_recording_done_pio_s1_begins_xfer;

  //vol_recording_done_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign vol_recording_done_pio_s1_in_a_read_cycle = cpu_data_master_granted_vol_recording_done_pio_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = vol_recording_done_pio_s1_in_a_read_cycle;

  //vol_recording_done_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign vol_recording_done_pio_s1_waits_for_write = vol_recording_done_pio_s1_in_a_write_cycle & 0;

  //vol_recording_done_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign vol_recording_done_pio_s1_in_a_write_cycle = cpu_data_master_granted_vol_recording_done_pio_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = vol_recording_done_pio_s1_in_a_write_cycle;

  assign wait_for_vol_recording_done_pio_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //vol_recording_done_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module vol_transfer_done_pio_s1_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_data_master_address_to_slave,
                                              cpu_data_master_latency_counter,
                                              cpu_data_master_read,
                                              cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register,
                                              cpu_data_master_write,
                                              cpu_data_master_writedata,
                                              reset_n,
                                              vol_transfer_done_pio_s1_readdata,

                                             // outputs:
                                              cpu_data_master_granted_vol_transfer_done_pio_s1,
                                              cpu_data_master_qualified_request_vol_transfer_done_pio_s1,
                                              cpu_data_master_read_data_valid_vol_transfer_done_pio_s1,
                                              cpu_data_master_requests_vol_transfer_done_pio_s1,
                                              d1_vol_transfer_done_pio_s1_end_xfer,
                                              vol_transfer_done_pio_s1_address,
                                              vol_transfer_done_pio_s1_chipselect,
                                              vol_transfer_done_pio_s1_readdata_from_sa,
                                              vol_transfer_done_pio_s1_reset_n,
                                              vol_transfer_done_pio_s1_write_n,
                                              vol_transfer_done_pio_s1_writedata
                                           )
;

  output           cpu_data_master_granted_vol_transfer_done_pio_s1;
  output           cpu_data_master_qualified_request_vol_transfer_done_pio_s1;
  output           cpu_data_master_read_data_valid_vol_transfer_done_pio_s1;
  output           cpu_data_master_requests_vol_transfer_done_pio_s1;
  output           d1_vol_transfer_done_pio_s1_end_xfer;
  output  [  1: 0] vol_transfer_done_pio_s1_address;
  output           vol_transfer_done_pio_s1_chipselect;
  output           vol_transfer_done_pio_s1_readdata_from_sa;
  output           vol_transfer_done_pio_s1_reset_n;
  output           vol_transfer_done_pio_s1_write_n;
  output           vol_transfer_done_pio_s1_writedata;
  input            clk;
  input   [ 30: 0] cpu_data_master_address_to_slave;
  input   [  1: 0] cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            vol_transfer_done_pio_s1_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_vol_transfer_done_pio_s1;
  wire             cpu_data_master_qualified_request_vol_transfer_done_pio_s1;
  wire             cpu_data_master_read_data_valid_vol_transfer_done_pio_s1;
  wire             cpu_data_master_requests_vol_transfer_done_pio_s1;
  wire             cpu_data_master_saved_grant_vol_transfer_done_pio_s1;
  reg              d1_reasons_to_wait;
  reg              d1_vol_transfer_done_pio_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 30: 0] shifted_address_to_vol_transfer_done_pio_s1_from_cpu_data_master;
  wire    [  1: 0] vol_transfer_done_pio_s1_address;
  wire             vol_transfer_done_pio_s1_allgrants;
  wire             vol_transfer_done_pio_s1_allow_new_arb_cycle;
  wire             vol_transfer_done_pio_s1_any_bursting_master_saved_grant;
  wire             vol_transfer_done_pio_s1_any_continuerequest;
  wire             vol_transfer_done_pio_s1_arb_counter_enable;
  reg     [  1: 0] vol_transfer_done_pio_s1_arb_share_counter;
  wire    [  1: 0] vol_transfer_done_pio_s1_arb_share_counter_next_value;
  wire    [  1: 0] vol_transfer_done_pio_s1_arb_share_set_values;
  wire             vol_transfer_done_pio_s1_beginbursttransfer_internal;
  wire             vol_transfer_done_pio_s1_begins_xfer;
  wire             vol_transfer_done_pio_s1_chipselect;
  wire             vol_transfer_done_pio_s1_end_xfer;
  wire             vol_transfer_done_pio_s1_firsttransfer;
  wire             vol_transfer_done_pio_s1_grant_vector;
  wire             vol_transfer_done_pio_s1_in_a_read_cycle;
  wire             vol_transfer_done_pio_s1_in_a_write_cycle;
  wire             vol_transfer_done_pio_s1_master_qreq_vector;
  wire             vol_transfer_done_pio_s1_non_bursting_master_requests;
  wire             vol_transfer_done_pio_s1_readdata_from_sa;
  reg              vol_transfer_done_pio_s1_reg_firsttransfer;
  wire             vol_transfer_done_pio_s1_reset_n;
  reg              vol_transfer_done_pio_s1_slavearbiterlockenable;
  wire             vol_transfer_done_pio_s1_slavearbiterlockenable2;
  wire             vol_transfer_done_pio_s1_unreg_firsttransfer;
  wire             vol_transfer_done_pio_s1_waits_for_read;
  wire             vol_transfer_done_pio_s1_waits_for_write;
  wire             vol_transfer_done_pio_s1_write_n;
  wire             vol_transfer_done_pio_s1_writedata;
  wire             wait_for_vol_transfer_done_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~vol_transfer_done_pio_s1_end_xfer;
    end


  assign vol_transfer_done_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_vol_transfer_done_pio_s1));
  //assign vol_transfer_done_pio_s1_readdata_from_sa = vol_transfer_done_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign vol_transfer_done_pio_s1_readdata_from_sa = vol_transfer_done_pio_s1_readdata;

  assign cpu_data_master_requests_vol_transfer_done_pio_s1 = ({cpu_data_master_address_to_slave[30 : 4] , 4'b0} == 31'h48112700) & (cpu_data_master_read | cpu_data_master_write);
  //vol_transfer_done_pio_s1_arb_share_counter set values, which is an e_mux
  assign vol_transfer_done_pio_s1_arb_share_set_values = 1;

  //vol_transfer_done_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign vol_transfer_done_pio_s1_non_bursting_master_requests = cpu_data_master_requests_vol_transfer_done_pio_s1;

  //vol_transfer_done_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign vol_transfer_done_pio_s1_any_bursting_master_saved_grant = 0;

  //vol_transfer_done_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign vol_transfer_done_pio_s1_arb_share_counter_next_value = vol_transfer_done_pio_s1_firsttransfer ? (vol_transfer_done_pio_s1_arb_share_set_values - 1) : |vol_transfer_done_pio_s1_arb_share_counter ? (vol_transfer_done_pio_s1_arb_share_counter - 1) : 0;

  //vol_transfer_done_pio_s1_allgrants all slave grants, which is an e_mux
  assign vol_transfer_done_pio_s1_allgrants = |vol_transfer_done_pio_s1_grant_vector;

  //vol_transfer_done_pio_s1_end_xfer assignment, which is an e_assign
  assign vol_transfer_done_pio_s1_end_xfer = ~(vol_transfer_done_pio_s1_waits_for_read | vol_transfer_done_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1 = vol_transfer_done_pio_s1_end_xfer & (~vol_transfer_done_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //vol_transfer_done_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign vol_transfer_done_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1 & vol_transfer_done_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1 & ~vol_transfer_done_pio_s1_non_bursting_master_requests);

  //vol_transfer_done_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_transfer_done_pio_s1_arb_share_counter <= 0;
      else if (vol_transfer_done_pio_s1_arb_counter_enable)
          vol_transfer_done_pio_s1_arb_share_counter <= vol_transfer_done_pio_s1_arb_share_counter_next_value;
    end


  //vol_transfer_done_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_transfer_done_pio_s1_slavearbiterlockenable <= 0;
      else if ((|vol_transfer_done_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1) | (end_xfer_arb_share_counter_term_vol_transfer_done_pio_s1 & ~vol_transfer_done_pio_s1_non_bursting_master_requests))
          vol_transfer_done_pio_s1_slavearbiterlockenable <= |vol_transfer_done_pio_s1_arb_share_counter_next_value;
    end


  //cpu/data_master vol_transfer_done_pio/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = vol_transfer_done_pio_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //vol_transfer_done_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign vol_transfer_done_pio_s1_slavearbiterlockenable2 = |vol_transfer_done_pio_s1_arb_share_counter_next_value;

  //cpu/data_master vol_transfer_done_pio/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = vol_transfer_done_pio_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //vol_transfer_done_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign vol_transfer_done_pio_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_vol_transfer_done_pio_s1 = cpu_data_master_requests_vol_transfer_done_pio_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_vol_transfer_done_pio_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_vol_transfer_done_pio_s1 = cpu_data_master_granted_vol_transfer_done_pio_s1 & cpu_data_master_read & ~vol_transfer_done_pio_s1_waits_for_read;

  //vol_transfer_done_pio_s1_writedata mux, which is an e_mux
  assign vol_transfer_done_pio_s1_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_vol_transfer_done_pio_s1 = cpu_data_master_qualified_request_vol_transfer_done_pio_s1;

  //cpu/data_master saved-grant vol_transfer_done_pio/s1, which is an e_assign
  assign cpu_data_master_saved_grant_vol_transfer_done_pio_s1 = cpu_data_master_requests_vol_transfer_done_pio_s1;

  //allow new arb cycle for vol_transfer_done_pio/s1, which is an e_assign
  assign vol_transfer_done_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign vol_transfer_done_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign vol_transfer_done_pio_s1_master_qreq_vector = 1;

  //vol_transfer_done_pio_s1_reset_n assignment, which is an e_assign
  assign vol_transfer_done_pio_s1_reset_n = reset_n;

  assign vol_transfer_done_pio_s1_chipselect = cpu_data_master_granted_vol_transfer_done_pio_s1;
  //vol_transfer_done_pio_s1_firsttransfer first transaction, which is an e_assign
  assign vol_transfer_done_pio_s1_firsttransfer = vol_transfer_done_pio_s1_begins_xfer ? vol_transfer_done_pio_s1_unreg_firsttransfer : vol_transfer_done_pio_s1_reg_firsttransfer;

  //vol_transfer_done_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign vol_transfer_done_pio_s1_unreg_firsttransfer = ~(vol_transfer_done_pio_s1_slavearbiterlockenable & vol_transfer_done_pio_s1_any_continuerequest);

  //vol_transfer_done_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          vol_transfer_done_pio_s1_reg_firsttransfer <= 1'b1;
      else if (vol_transfer_done_pio_s1_begins_xfer)
          vol_transfer_done_pio_s1_reg_firsttransfer <= vol_transfer_done_pio_s1_unreg_firsttransfer;
    end


  //vol_transfer_done_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign vol_transfer_done_pio_s1_beginbursttransfer_internal = vol_transfer_done_pio_s1_begins_xfer;

  //~vol_transfer_done_pio_s1_write_n assignment, which is an e_mux
  assign vol_transfer_done_pio_s1_write_n = ~(cpu_data_master_granted_vol_transfer_done_pio_s1 & cpu_data_master_write);

  assign shifted_address_to_vol_transfer_done_pio_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //vol_transfer_done_pio_s1_address mux, which is an e_mux
  assign vol_transfer_done_pio_s1_address = shifted_address_to_vol_transfer_done_pio_s1_from_cpu_data_master >> 2;

  //d1_vol_transfer_done_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_vol_transfer_done_pio_s1_end_xfer <= 1;
      else 
        d1_vol_transfer_done_pio_s1_end_xfer <= vol_transfer_done_pio_s1_end_xfer;
    end


  //vol_transfer_done_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign vol_transfer_done_pio_s1_waits_for_read = vol_transfer_done_pio_s1_in_a_read_cycle & vol_transfer_done_pio_s1_begins_xfer;

  //vol_transfer_done_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign vol_transfer_done_pio_s1_in_a_read_cycle = cpu_data_master_granted_vol_transfer_done_pio_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = vol_transfer_done_pio_s1_in_a_read_cycle;

  //vol_transfer_done_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign vol_transfer_done_pio_s1_waits_for_write = vol_transfer_done_pio_s1_in_a_write_cycle & 0;

  //vol_transfer_done_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign vol_transfer_done_pio_s1_in_a_write_cycle = cpu_data_master_granted_vol_transfer_done_pio_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = vol_transfer_done_pio_s1_in_a_write_cycle;

  assign wait_for_vol_transfer_done_pio_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //vol_transfer_done_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_reset_ddr2_phy_clk_out_domain_synch_module (
                                                                // inputs:
                                                                 clk,
                                                                 data_in,
                                                                 reset_n,

                                                                // outputs:
                                                                 data_out
                                                              )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC_reset_pll_sys_clk_domain_synch_module (
                                                           // inputs:
                                                            clk,
                                                            data_in,
                                                            reset_n,

                                                           // outputs:
                                                            data_out
                                                         )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module SS_OCT_SOPC (
                     // 1) global signals:
                      clk_50,
                      ddr2_aux_full_rate_clk_out,
                      ddr2_aux_half_rate_clk_out,
                      ddr2_phy_clk_out,
                      pll_sys_clk,
                      reset_n,

                     // the_ddr2
                      aux_scan_clk_from_the_ddr2,
                      aux_scan_clk_reset_n_from_the_ddr2,
                      dll_reference_clk_from_the_ddr2,
                      dqs_delay_ctrl_export_from_the_ddr2,
                      global_reset_n_to_the_ddr2,
                      local_init_done_from_the_ddr2,
                      local_refresh_ack_from_the_ddr2,
                      local_wdata_req_from_the_ddr2,
                      mem_addr_from_the_ddr2,
                      mem_ba_from_the_ddr2,
                      mem_cas_n_from_the_ddr2,
                      mem_cke_from_the_ddr2,
                      mem_clk_n_to_and_from_the_ddr2,
                      mem_clk_to_and_from_the_ddr2,
                      mem_cs_n_from_the_ddr2,
                      mem_dm_from_the_ddr2,
                      mem_dq_to_and_from_the_ddr2,
                      mem_dqs_to_and_from_the_ddr2,
                      mem_dqsn_to_and_from_the_ddr2,
                      mem_odt_from_the_ddr2,
                      mem_ras_n_from_the_ddr2,
                      mem_we_n_from_the_ddr2,
                      oct_ctl_rs_value_to_the_ddr2,
                      oct_ctl_rt_value_to_the_ddr2,
                      reset_phy_clk_n_from_the_ddr2,

                     // the_flash_tristate_bridge_avalon_slave
                      flash_tristate_bridge_address,
                      flash_tristate_bridge_data,
                      flash_tristate_bridge_readn,
                      flash_tristate_bridge_writen,
                      select_n_to_the_ext_flash,

                     // the_master_read
                      control_done_from_the_master_read,
                      control_early_done_from_the_master_read,
                      control_fixed_location_to_the_master_read,
                      control_go_to_the_master_read,
                      control_read_base_to_the_master_read,
                      control_read_length_to_the_master_read,
                      user_buffer_output_data_from_the_master_read,
                      user_data_available_from_the_master_read,
                      user_read_buffer_to_the_master_read,

                     // the_master_write
                      control_done_from_the_master_write,
                      control_fixed_location_to_the_master_write,
                      control_go_to_the_master_write,
                      control_write_base_to_the_master_write,
                      control_write_length_to_the_master_write,
                      user_buffer_full_from_the_master_write,
                      user_buffer_input_data_to_the_master_write,
                      user_write_buffer_to_the_master_write,

                     // the_tse_mac
                      led_an_from_the_tse_mac,
                      led_char_err_from_the_tse_mac,
                      led_col_from_the_tse_mac,
                      led_crs_from_the_tse_mac,
                      led_disp_err_from_the_tse_mac,
                      led_link_from_the_tse_mac,
                      mdc_from_the_tse_mac,
                      mdio_in_to_the_tse_mac,
                      mdio_oen_from_the_tse_mac,
                      mdio_out_from_the_tse_mac,
                      ref_clk_to_the_tse_mac,
                      rxp_to_the_tse_mac,
                      txp_from_the_tse_mac,

                     // the_vol_recording_done_pio
                      in_port_to_the_vol_recording_done_pio,

                     // the_vol_transfer_done_pio
                      out_port_from_the_vol_transfer_done_pio
                   )
;

  output           aux_scan_clk_from_the_ddr2;
  output           aux_scan_clk_reset_n_from_the_ddr2;
  output           control_done_from_the_master_read;
  output           control_done_from_the_master_write;
  output           control_early_done_from_the_master_read;
  output           ddr2_aux_full_rate_clk_out;
  output           ddr2_aux_half_rate_clk_out;
  output           ddr2_phy_clk_out;
  output           dll_reference_clk_from_the_ddr2;
  output  [  5: 0] dqs_delay_ctrl_export_from_the_ddr2;
  output  [ 25: 0] flash_tristate_bridge_address;
  inout   [ 15: 0] flash_tristate_bridge_data;
  output           flash_tristate_bridge_readn;
  output           flash_tristate_bridge_writen;
  output           led_an_from_the_tse_mac;
  output           led_char_err_from_the_tse_mac;
  output           led_col_from_the_tse_mac;
  output           led_crs_from_the_tse_mac;
  output           led_disp_err_from_the_tse_mac;
  output           led_link_from_the_tse_mac;
  output           local_init_done_from_the_ddr2;
  output           local_refresh_ack_from_the_ddr2;
  output           local_wdata_req_from_the_ddr2;
  output           mdc_from_the_tse_mac;
  output           mdio_oen_from_the_tse_mac;
  output           mdio_out_from_the_tse_mac;
  output  [ 13: 0] mem_addr_from_the_ddr2;
  output  [  2: 0] mem_ba_from_the_ddr2;
  output           mem_cas_n_from_the_ddr2;
  output           mem_cke_from_the_ddr2;
  inout   [  1: 0] mem_clk_n_to_and_from_the_ddr2;
  inout   [  1: 0] mem_clk_to_and_from_the_ddr2;
  output           mem_cs_n_from_the_ddr2;
  output  [  7: 0] mem_dm_from_the_ddr2;
  inout   [ 63: 0] mem_dq_to_and_from_the_ddr2;
  inout   [  7: 0] mem_dqs_to_and_from_the_ddr2;
  inout   [  7: 0] mem_dqsn_to_and_from_the_ddr2;
  output           mem_odt_from_the_ddr2;
  output           mem_ras_n_from_the_ddr2;
  output           mem_we_n_from_the_ddr2;
  output           out_port_from_the_vol_transfer_done_pio;
  output           pll_sys_clk;
  output           reset_phy_clk_n_from_the_ddr2;
  output           select_n_to_the_ext_flash;
  output           txp_from_the_tse_mac;
  output           user_buffer_full_from_the_master_write;
  output  [255: 0] user_buffer_output_data_from_the_master_read;
  output           user_data_available_from_the_master_read;
  input            clk_50;
  input            control_fixed_location_to_the_master_read;
  input            control_fixed_location_to_the_master_write;
  input            control_go_to_the_master_read;
  input            control_go_to_the_master_write;
  input   [ 29: 0] control_read_base_to_the_master_read;
  input   [ 29: 0] control_read_length_to_the_master_read;
  input   [ 29: 0] control_write_base_to_the_master_write;
  input   [ 29: 0] control_write_length_to_the_master_write;
  input            global_reset_n_to_the_ddr2;
  input            in_port_to_the_vol_recording_done_pio;
  input            mdio_in_to_the_tse_mac;
  input   [ 13: 0] oct_ctl_rs_value_to_the_ddr2;
  input   [ 13: 0] oct_ctl_rt_value_to_the_ddr2;
  input            ref_clk_to_the_tse_mac;
  input            reset_n;
  input            rxp_to_the_tse_mac;
  input   [255: 0] user_buffer_input_data_to_the_master_write;
  input            user_read_buffer_to_the_master_read;
  input            user_write_buffer_to_the_master_write;

  wire    [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address;
  wire    [ 29: 0] SS_OCT_SOPC_burst_0_downstream_address_to_slave;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_downstream_arbitrationshare;
  wire    [  2: 0] SS_OCT_SOPC_burst_0_downstream_burstcount;
  wire    [ 31: 0] SS_OCT_SOPC_burst_0_downstream_byteenable;
  wire             SS_OCT_SOPC_burst_0_downstream_debugaccess;
  wire             SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_latency_counter;
  wire    [ 29: 0] SS_OCT_SOPC_burst_0_downstream_nativeaddress;
  wire             SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_read;
  wire             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register;
  wire    [255: 0] SS_OCT_SOPC_burst_0_downstream_readdata;
  wire             SS_OCT_SOPC_burst_0_downstream_readdatavalid;
  wire             SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1;
  wire             SS_OCT_SOPC_burst_0_downstream_reset_n;
  wire             SS_OCT_SOPC_burst_0_downstream_waitrequest;
  wire             SS_OCT_SOPC_burst_0_downstream_write;
  wire    [255: 0] SS_OCT_SOPC_burst_0_downstream_writedata;
  wire    [ 29: 0] SS_OCT_SOPC_burst_0_upstream_address;
  wire    [  3: 0] SS_OCT_SOPC_burst_0_upstream_burstcount;
  wire    [ 34: 0] SS_OCT_SOPC_burst_0_upstream_byteaddress;
  wire    [ 31: 0] SS_OCT_SOPC_burst_0_upstream_byteenable;
  wire             SS_OCT_SOPC_burst_0_upstream_debugaccess;
  wire             SS_OCT_SOPC_burst_0_upstream_read;
  wire    [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata;
  wire    [255: 0] SS_OCT_SOPC_burst_0_upstream_readdata_from_sa;
  wire             SS_OCT_SOPC_burst_0_upstream_readdatavalid;
  wire             SS_OCT_SOPC_burst_0_upstream_waitrequest;
  wire             SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa;
  wire             SS_OCT_SOPC_burst_0_upstream_write;
  wire    [255: 0] SS_OCT_SOPC_burst_0_upstream_writedata;
  wire    [  3: 0] SS_OCT_SOPC_clock_0_in_address;
  wire    [  1: 0] SS_OCT_SOPC_clock_0_in_byteenable;
  wire             SS_OCT_SOPC_clock_0_in_endofpacket;
  wire             SS_OCT_SOPC_clock_0_in_endofpacket_from_sa;
  wire    [  2: 0] SS_OCT_SOPC_clock_0_in_nativeaddress;
  wire             SS_OCT_SOPC_clock_0_in_read;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_in_readdata_from_sa;
  wire             SS_OCT_SOPC_clock_0_in_reset_n;
  wire             SS_OCT_SOPC_clock_0_in_waitrequest;
  wire             SS_OCT_SOPC_clock_0_in_waitrequest_from_sa;
  wire             SS_OCT_SOPC_clock_0_in_write;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_in_writedata;
  wire    [  3: 0] SS_OCT_SOPC_clock_0_out_address;
  wire    [  3: 0] SS_OCT_SOPC_clock_0_out_address_to_slave;
  wire    [  1: 0] SS_OCT_SOPC_clock_0_out_byteenable;
  wire             SS_OCT_SOPC_clock_0_out_endofpacket;
  wire             SS_OCT_SOPC_clock_0_out_granted_pll_s1;
  wire    [  2: 0] SS_OCT_SOPC_clock_0_out_nativeaddress;
  wire             SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_read;
  wire             SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_out_readdata;
  wire             SS_OCT_SOPC_clock_0_out_requests_pll_s1;
  wire             SS_OCT_SOPC_clock_0_out_reset_n;
  wire             SS_OCT_SOPC_clock_0_out_waitrequest;
  wire             SS_OCT_SOPC_clock_0_out_write;
  wire    [ 15: 0] SS_OCT_SOPC_clock_0_out_writedata;
  wire             aux_scan_clk_from_the_ddr2;
  wire             aux_scan_clk_reset_n_from_the_ddr2;
  wire             clk_50_reset_n;
  wire    [ 29: 0] clock_crossing_ddr2_cpu_m1_address;
  wire    [ 29: 0] clock_crossing_ddr2_cpu_m1_address_to_slave;
  wire    [  3: 0] clock_crossing_ddr2_cpu_m1_byteenable;
  wire             clock_crossing_ddr2_cpu_m1_endofpacket;
  wire             clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_latency_counter;
  wire    [ 27: 0] clock_crossing_ddr2_cpu_m1_nativeaddress;
  wire             clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_read;
  wire             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_m1_readdata;
  wire             clock_crossing_ddr2_cpu_m1_readdatavalid;
  wire             clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1;
  wire             clock_crossing_ddr2_cpu_m1_reset_n;
  wire             clock_crossing_ddr2_cpu_m1_waitrequest;
  wire             clock_crossing_ddr2_cpu_m1_write;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_m1_writedata;
  wire    [ 27: 0] clock_crossing_ddr2_cpu_s1_address;
  wire    [  3: 0] clock_crossing_ddr2_cpu_s1_byteenable;
  wire             clock_crossing_ddr2_cpu_s1_endofpacket;
  wire             clock_crossing_ddr2_cpu_s1_endofpacket_from_sa;
  wire    [ 27: 0] clock_crossing_ddr2_cpu_s1_nativeaddress;
  wire             clock_crossing_ddr2_cpu_s1_read;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_s1_readdata_from_sa;
  wire             clock_crossing_ddr2_cpu_s1_readdatavalid;
  wire             clock_crossing_ddr2_cpu_s1_reset_n;
  wire             clock_crossing_ddr2_cpu_s1_waitrequest;
  wire             clock_crossing_ddr2_cpu_s1_waitrequest_from_sa;
  wire             clock_crossing_ddr2_cpu_s1_write;
  wire    [ 31: 0] clock_crossing_ddr2_cpu_s1_writedata;
  wire    [ 29: 0] clock_crossing_master_ddr2_m1_address;
  wire    [ 29: 0] clock_crossing_master_ddr2_m1_address_to_slave;
  wire    [  3: 0] clock_crossing_master_ddr2_m1_burstcount;
  wire    [ 31: 0] clock_crossing_master_ddr2_m1_byteenable;
  wire             clock_crossing_master_ddr2_m1_endofpacket;
  wire             clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_latency_counter;
  wire    [ 24: 0] clock_crossing_master_ddr2_m1_nativeaddress;
  wire             clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_read;
  wire             clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register;
  wire    [255: 0] clock_crossing_master_ddr2_m1_readdata;
  wire             clock_crossing_master_ddr2_m1_readdatavalid;
  wire             clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream;
  wire             clock_crossing_master_ddr2_m1_reset_n;
  wire             clock_crossing_master_ddr2_m1_waitrequest;
  wire             clock_crossing_master_ddr2_m1_write;
  wire    [255: 0] clock_crossing_master_ddr2_m1_writedata;
  wire    [ 24: 0] clock_crossing_master_ddr2_s1_address;
  wire    [  3: 0] clock_crossing_master_ddr2_s1_burstcount;
  wire    [ 31: 0] clock_crossing_master_ddr2_s1_byteenable;
  wire             clock_crossing_master_ddr2_s1_endofpacket;
  wire             clock_crossing_master_ddr2_s1_endofpacket_from_sa;
  wire    [ 24: 0] clock_crossing_master_ddr2_s1_nativeaddress;
  wire             clock_crossing_master_ddr2_s1_read;
  wire    [255: 0] clock_crossing_master_ddr2_s1_readdata;
  wire    [255: 0] clock_crossing_master_ddr2_s1_readdata_from_sa;
  wire             clock_crossing_master_ddr2_s1_readdatavalid;
  wire             clock_crossing_master_ddr2_s1_reset_n;
  wire             clock_crossing_master_ddr2_s1_waitrequest;
  wire             clock_crossing_master_ddr2_s1_waitrequest_from_sa;
  wire             clock_crossing_master_ddr2_s1_write;
  wire    [255: 0] clock_crossing_master_ddr2_s1_writedata;
  wire             control_done_from_the_master_read;
  wire             control_done_from_the_master_write;
  wire             control_early_done_from_the_master_read;
  wire    [ 30: 0] cpu_data_master_address;
  wire    [ 30: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire    [  1: 0] cpu_data_master_byteenable_ext_flash_s1;
  wire    [  1: 0] cpu_data_master_dbs_address;
  wire    [ 15: 0] cpu_data_master_dbs_write_16;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_granted_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_granted_descriptor_memory_s1;
  wire             cpu_data_master_granted_ext_flash_s1;
  wire             cpu_data_master_granted_high_res_timer_s1;
  wire             cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_granted_onchip_memory_s1;
  wire             cpu_data_master_granted_packet_memory_s1;
  wire             cpu_data_master_granted_sgdma_rx_csr;
  wire             cpu_data_master_granted_sgdma_tx_csr;
  wire             cpu_data_master_granted_sys_timer_s1;
  wire             cpu_data_master_granted_sysid_control_slave;
  wire             cpu_data_master_granted_tse_mac_control_port;
  wire             cpu_data_master_granted_vol_recording_done_pio_s1;
  wire             cpu_data_master_granted_vol_transfer_done_pio_s1;
  wire    [ 31: 0] cpu_data_master_irq;
  wire    [  1: 0] cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_descriptor_memory_s1;
  wire             cpu_data_master_qualified_request_ext_flash_s1;
  wire             cpu_data_master_qualified_request_high_res_timer_s1;
  wire             cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_qualified_request_onchip_memory_s1;
  wire             cpu_data_master_qualified_request_packet_memory_s1;
  wire             cpu_data_master_qualified_request_sgdma_rx_csr;
  wire             cpu_data_master_qualified_request_sgdma_tx_csr;
  wire             cpu_data_master_qualified_request_sys_timer_s1;
  wire             cpu_data_master_qualified_request_sysid_control_slave;
  wire             cpu_data_master_qualified_request_tse_mac_control_port;
  wire             cpu_data_master_qualified_request_vol_recording_done_pio_s1;
  wire             cpu_data_master_qualified_request_vol_transfer_done_pio_s1;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1;
  wire             cpu_data_master_read_data_valid_ext_flash_s1;
  wire             cpu_data_master_read_data_valid_high_res_timer_s1;
  wire             cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_read_data_valid_onchip_memory_s1;
  wire             cpu_data_master_read_data_valid_packet_memory_s1;
  wire             cpu_data_master_read_data_valid_sgdma_rx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_tx_csr;
  wire             cpu_data_master_read_data_valid_sys_timer_s1;
  wire             cpu_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_data_master_read_data_valid_tse_mac_control_port;
  wire             cpu_data_master_read_data_valid_vol_recording_done_pio_s1;
  wire             cpu_data_master_read_data_valid_vol_transfer_done_pio_s1;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_SS_OCT_SOPC_clock_0_in;
  wire             cpu_data_master_requests_clock_crossing_ddr2_cpu_s1;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_descriptor_memory_s1;
  wire             cpu_data_master_requests_ext_flash_s1;
  wire             cpu_data_master_requests_high_res_timer_s1;
  wire             cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  wire             cpu_data_master_requests_onchip_memory_s1;
  wire             cpu_data_master_requests_packet_memory_s1;
  wire             cpu_data_master_requests_sgdma_rx_csr;
  wire             cpu_data_master_requests_sgdma_tx_csr;
  wire             cpu_data_master_requests_sys_timer_s1;
  wire             cpu_data_master_requests_sysid_control_slave;
  wire             cpu_data_master_requests_tse_mac_control_port;
  wire             cpu_data_master_requests_vol_recording_done_pio_s1;
  wire             cpu_data_master_requests_vol_transfer_done_pio_s1;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 30: 0] cpu_instruction_master_address;
  wire    [ 30: 0] cpu_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_instruction_master_dbs_address;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_granted_descriptor_memory_s1;
  wire             cpu_instruction_master_granted_ext_flash_s1;
  wire             cpu_instruction_master_granted_onchip_memory_s1;
  wire    [  1: 0] cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_descriptor_memory_s1;
  wire             cpu_instruction_master_qualified_request_ext_flash_s1;
  wire             cpu_instruction_master_qualified_request_onchip_memory_s1;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_descriptor_memory_s1;
  wire             cpu_instruction_master_read_data_valid_ext_flash_s1;
  wire             cpu_instruction_master_read_data_valid_onchip_memory_s1;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_descriptor_memory_s1;
  wire             cpu_instruction_master_requests_ext_flash_s1;
  wire             cpu_instruction_master_requests_onchip_memory_s1;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire             d1_SS_OCT_SOPC_burst_0_upstream_end_xfer;
  wire             d1_SS_OCT_SOPC_clock_0_in_end_xfer;
  wire             d1_clock_crossing_ddr2_cpu_s1_end_xfer;
  wire             d1_clock_crossing_master_ddr2_s1_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_ddr2_s1_end_xfer;
  wire             d1_descriptor_memory_s1_end_xfer;
  wire             d1_flash_tristate_bridge_avalon_slave_end_xfer;
  wire             d1_high_res_timer_s1_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_onchip_memory_s1_end_xfer;
  wire             d1_packet_memory_s1_end_xfer;
  wire             d1_packet_memory_s2_end_xfer;
  wire             d1_pipeline_bridge_ddr2_s1_end_xfer;
  wire             d1_pll_s1_end_xfer;
  wire             d1_sgdma_rx_csr_end_xfer;
  wire             d1_sgdma_tx_csr_end_xfer;
  wire             d1_sys_timer_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_tse_mac_control_port_end_xfer;
  wire             d1_vol_recording_done_pio_s1_end_xfer;
  wire             d1_vol_transfer_done_pio_s1_end_xfer;
  wire             ddr2_aux_full_rate_clk_out;
  wire             ddr2_aux_half_rate_clk_out;
  wire             ddr2_phy_clk_out;
  wire             ddr2_phy_clk_out_reset_n;
  wire    [ 24: 0] ddr2_s1_address;
  wire             ddr2_s1_beginbursttransfer;
  wire    [  2: 0] ddr2_s1_burstcount;
  wire    [ 31: 0] ddr2_s1_byteenable;
  wire             ddr2_s1_read;
  wire    [255: 0] ddr2_s1_readdata;
  wire    [255: 0] ddr2_s1_readdata_from_sa;
  wire             ddr2_s1_readdatavalid;
  wire             ddr2_s1_resetrequest_n;
  wire             ddr2_s1_resetrequest_n_from_sa;
  wire             ddr2_s1_waitrequest_n;
  wire             ddr2_s1_waitrequest_n_from_sa;
  wire             ddr2_s1_write;
  wire    [255: 0] ddr2_s1_writedata;
  wire    [  8: 0] descriptor_memory_s1_address;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire             descriptor_memory_s1_clken;
  wire    [ 31: 0] descriptor_memory_s1_readdata;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  wire             dll_reference_clk_from_the_ddr2;
  wire    [  5: 0] dqs_delay_ctrl_export_from_the_ddr2;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire    [ 25: 0] flash_tristate_bridge_address;
  wire    [ 15: 0] flash_tristate_bridge_data;
  wire             flash_tristate_bridge_readn;
  wire             flash_tristate_bridge_writen;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_irq;
  wire             high_res_timer_s1_irq_from_sa;
  wire    [ 15: 0] high_res_timer_s1_readdata;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  wire             high_res_timer_s1_reset_n;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire    [ 15: 0] incoming_flash_tristate_bridge_data;
  wire    [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             led_an_from_the_tse_mac;
  wire             led_char_err_from_the_tse_mac;
  wire             led_col_from_the_tse_mac;
  wire             led_crs_from_the_tse_mac;
  wire             led_disp_err_from_the_tse_mac;
  wire             led_link_from_the_tse_mac;
  wire             local_init_done_from_the_ddr2;
  wire             local_refresh_ack_from_the_ddr2;
  wire             local_wdata_req_from_the_ddr2;
  wire    [ 29: 0] master_read_avalon_master_address;
  wire    [ 29: 0] master_read_avalon_master_address_to_slave;
  wire    [  3: 0] master_read_avalon_master_burstcount;
  wire    [ 31: 0] master_read_avalon_master_byteenable;
  wire             master_read_avalon_master_read;
  wire    [255: 0] master_read_avalon_master_readdata;
  wire             master_read_avalon_master_readdatavalid;
  wire             master_read_avalon_master_reset;
  wire             master_read_avalon_master_waitrequest;
  wire             master_read_granted_clock_crossing_master_ddr2_s1;
  wire             master_read_latency_counter;
  wire             master_read_qualified_request_clock_crossing_master_ddr2_s1;
  wire             master_read_read_data_valid_clock_crossing_master_ddr2_s1;
  wire             master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register;
  wire             master_read_requests_clock_crossing_master_ddr2_s1;
  wire    [ 29: 0] master_write_avalon_master_address;
  wire    [ 29: 0] master_write_avalon_master_address_to_slave;
  wire    [  3: 0] master_write_avalon_master_burstcount;
  wire    [ 31: 0] master_write_avalon_master_byteenable;
  wire             master_write_avalon_master_reset;
  wire             master_write_avalon_master_waitrequest;
  wire             master_write_avalon_master_write;
  wire    [255: 0] master_write_avalon_master_writedata;
  wire             master_write_granted_clock_crossing_master_ddr2_s1;
  wire             master_write_qualified_request_clock_crossing_master_ddr2_s1;
  wire             master_write_requests_clock_crossing_master_ddr2_s1;
  wire             mdc_from_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 13: 0] mem_addr_from_the_ddr2;
  wire    [  2: 0] mem_ba_from_the_ddr2;
  wire             mem_cas_n_from_the_ddr2;
  wire             mem_cke_from_the_ddr2;
  wire    [  1: 0] mem_clk_n_to_and_from_the_ddr2;
  wire    [  1: 0] mem_clk_to_and_from_the_ddr2;
  wire             mem_cs_n_from_the_ddr2;
  wire    [  7: 0] mem_dm_from_the_ddr2;
  wire    [ 63: 0] mem_dq_to_and_from_the_ddr2;
  wire    [  7: 0] mem_dqs_to_and_from_the_ddr2;
  wire    [  7: 0] mem_dqsn_to_and_from_the_ddr2;
  wire             mem_odt_from_the_ddr2;
  wire             mem_ras_n_from_the_ddr2;
  wire             mem_we_n_from_the_ddr2;
  wire    [ 16: 0] onchip_memory_s1_address;
  wire    [  3: 0] onchip_memory_s1_byteenable;
  wire             onchip_memory_s1_chipselect;
  wire             onchip_memory_s1_clken;
  wire    [ 31: 0] onchip_memory_s1_readdata;
  wire    [ 31: 0] onchip_memory_s1_readdata_from_sa;
  wire             onchip_memory_s1_write;
  wire    [ 31: 0] onchip_memory_s1_writedata;
  wire             out_clk_ddr2_aux_full_rate_clk;
  wire             out_clk_ddr2_aux_half_rate_clk;
  wire             out_clk_ddr2_phy_clk;
  wire             out_clk_pll_c0;
  wire             out_port_from_the_vol_transfer_done_pio;
  wire    [ 13: 0] packet_memory_s1_address;
  wire    [  3: 0] packet_memory_s1_byteenable;
  wire             packet_memory_s1_chipselect;
  wire             packet_memory_s1_clken;
  wire    [ 31: 0] packet_memory_s1_readdata;
  wire    [ 31: 0] packet_memory_s1_readdata_from_sa;
  wire             packet_memory_s1_write;
  wire    [ 31: 0] packet_memory_s1_writedata;
  wire    [ 13: 0] packet_memory_s2_address;
  wire    [  3: 0] packet_memory_s2_byteenable;
  wire             packet_memory_s2_chipselect;
  wire             packet_memory_s2_clken;
  wire    [ 31: 0] packet_memory_s2_readdata;
  wire    [ 31: 0] packet_memory_s2_readdata_from_sa;
  wire             packet_memory_s2_write;
  wire    [ 31: 0] packet_memory_s2_writedata;
  wire    [ 29: 0] pipeline_bridge_ddr2_m1_address;
  wire    [ 29: 0] pipeline_bridge_ddr2_m1_address_to_slave;
  wire             pipeline_bridge_ddr2_m1_burstcount;
  wire    [  3: 0] pipeline_bridge_ddr2_m1_byteenable;
  wire             pipeline_bridge_ddr2_m1_chipselect;
  wire             pipeline_bridge_ddr2_m1_debugaccess;
  wire             pipeline_bridge_ddr2_m1_endofpacket;
  wire             pipeline_bridge_ddr2_m1_granted_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_latency_counter;
  wire             pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_read;
  wire             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register;
  wire    [ 31: 0] pipeline_bridge_ddr2_m1_readdata;
  wire             pipeline_bridge_ddr2_m1_readdatavalid;
  wire             pipeline_bridge_ddr2_m1_requests_ddr2_s1;
  wire             pipeline_bridge_ddr2_m1_waitrequest;
  wire             pipeline_bridge_ddr2_m1_write;
  wire    [ 31: 0] pipeline_bridge_ddr2_m1_writedata;
  wire    [ 27: 0] pipeline_bridge_ddr2_s1_address;
  wire             pipeline_bridge_ddr2_s1_arbiterlock;
  wire             pipeline_bridge_ddr2_s1_arbiterlock2;
  wire             pipeline_bridge_ddr2_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_ddr2_s1_byteenable;
  wire             pipeline_bridge_ddr2_s1_chipselect;
  wire             pipeline_bridge_ddr2_s1_debugaccess;
  wire             pipeline_bridge_ddr2_s1_endofpacket;
  wire             pipeline_bridge_ddr2_s1_endofpacket_from_sa;
  wire    [ 27: 0] pipeline_bridge_ddr2_s1_nativeaddress;
  wire             pipeline_bridge_ddr2_s1_read;
  wire    [ 31: 0] pipeline_bridge_ddr2_s1_readdata;
  wire    [ 31: 0] pipeline_bridge_ddr2_s1_readdata_from_sa;
  wire             pipeline_bridge_ddr2_s1_readdatavalid;
  wire             pipeline_bridge_ddr2_s1_reset_n;
  wire             pipeline_bridge_ddr2_s1_waitrequest;
  wire             pipeline_bridge_ddr2_s1_waitrequest_from_sa;
  wire             pipeline_bridge_ddr2_s1_write;
  wire    [ 31: 0] pipeline_bridge_ddr2_s1_writedata;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_chipselect;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest;
  wire             pll_s1_resetrequest_from_sa;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             pll_sys_clk;
  wire             pll_sys_clk_reset_n;
  wire             reset_n_sources;
  wire             reset_phy_clk_n_from_the_ddr2;
  wire             select_n_to_the_ext_flash;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_irq;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  wire             sgdma_rx_csr_reset_n;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_latency_counter;
  wire             sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_waitrequest;
  wire             sgdma_rx_descriptor_write_write;
  wire    [ 31: 0] sgdma_rx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  3: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  wire    [ 31: 0] sgdma_rx_m_write_address;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  wire    [  3: 0] sgdma_rx_m_write_byteenable;
  wire             sgdma_rx_m_write_granted_onchip_memory_s1;
  wire             sgdma_rx_m_write_granted_packet_memory_s2;
  wire             sgdma_rx_m_write_qualified_request_onchip_memory_s1;
  wire             sgdma_rx_m_write_qualified_request_packet_memory_s2;
  wire             sgdma_rx_m_write_requests_onchip_memory_s1;
  wire             sgdma_rx_m_write_requests_packet_memory_s2;
  wire             sgdma_rx_m_write_waitrequest;
  wire             sgdma_rx_m_write_write;
  wire    [ 31: 0] sgdma_rx_m_write_writedata;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_irq;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  wire             sgdma_tx_csr_reset_n;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_latency_counter;
  wire             sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_waitrequest;
  wire             sgdma_tx_descriptor_write_write;
  wire    [ 31: 0] sgdma_tx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_tx_m_read_address;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_granted_onchip_memory_s1;
  wire             sgdma_tx_m_read_granted_packet_memory_s2;
  wire             sgdma_tx_m_read_latency_counter;
  wire             sgdma_tx_m_read_qualified_request_onchip_memory_s1;
  wire             sgdma_tx_m_read_qualified_request_packet_memory_s2;
  wire             sgdma_tx_m_read_read;
  wire             sgdma_tx_m_read_read_data_valid_onchip_memory_s1;
  wire             sgdma_tx_m_read_read_data_valid_packet_memory_s2;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_requests_onchip_memory_s1;
  wire             sgdma_tx_m_read_requests_packet_memory_s2;
  wire             sgdma_tx_m_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_out_data;
  wire    [  1: 0] sgdma_tx_out_empty;
  wire             sgdma_tx_out_endofpacket;
  wire             sgdma_tx_out_error;
  wire             sgdma_tx_out_ready;
  wire             sgdma_tx_out_startofpacket;
  wire             sgdma_tx_out_valid;
  wire    [  2: 0] sys_timer_s1_address;
  wire             sys_timer_s1_chipselect;
  wire             sys_timer_s1_irq;
  wire             sys_timer_s1_irq_from_sa;
  wire    [ 15: 0] sys_timer_s1_readdata;
  wire    [ 15: 0] sys_timer_s1_readdata_from_sa;
  wire             sys_timer_s1_reset_n;
  wire             sys_timer_s1_write_n;
  wire    [ 15: 0] sys_timer_s1_writedata;
  wire             sysid_control_slave_address;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  wire             tse_mac_control_port_reset;
  wire             tse_mac_control_port_waitrequest;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire    [ 31: 0] tse_mac_receive_data;
  wire    [  1: 0] tse_mac_receive_empty;
  wire             tse_mac_receive_endofpacket;
  wire    [  5: 0] tse_mac_receive_error;
  wire             tse_mac_receive_ready;
  wire             tse_mac_receive_startofpacket;
  wire             tse_mac_receive_valid;
  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  wire             txp_from_the_tse_mac;
  wire             user_buffer_full_from_the_master_write;
  wire    [255: 0] user_buffer_output_data_from_the_master_read;
  wire             user_data_available_from_the_master_read;
  wire    [  1: 0] vol_recording_done_pio_s1_address;
  wire             vol_recording_done_pio_s1_readdata;
  wire             vol_recording_done_pio_s1_readdata_from_sa;
  wire             vol_recording_done_pio_s1_reset_n;
  wire    [  1: 0] vol_transfer_done_pio_s1_address;
  wire             vol_transfer_done_pio_s1_chipselect;
  wire             vol_transfer_done_pio_s1_readdata;
  wire             vol_transfer_done_pio_s1_readdata_from_sa;
  wire             vol_transfer_done_pio_s1_reset_n;
  wire             vol_transfer_done_pio_s1_write_n;
  wire             vol_transfer_done_pio_s1_writedata;
  SS_OCT_SOPC_burst_0_upstream_arbitrator the_SS_OCT_SOPC_burst_0_upstream
    (
      .SS_OCT_SOPC_burst_0_upstream_address                                                      (SS_OCT_SOPC_burst_0_upstream_address),
      .SS_OCT_SOPC_burst_0_upstream_burstcount                                                   (SS_OCT_SOPC_burst_0_upstream_burstcount),
      .SS_OCT_SOPC_burst_0_upstream_byteaddress                                                  (SS_OCT_SOPC_burst_0_upstream_byteaddress),
      .SS_OCT_SOPC_burst_0_upstream_byteenable                                                   (SS_OCT_SOPC_burst_0_upstream_byteenable),
      .SS_OCT_SOPC_burst_0_upstream_debugaccess                                                  (SS_OCT_SOPC_burst_0_upstream_debugaccess),
      .SS_OCT_SOPC_burst_0_upstream_read                                                         (SS_OCT_SOPC_burst_0_upstream_read),
      .SS_OCT_SOPC_burst_0_upstream_readdata                                                     (SS_OCT_SOPC_burst_0_upstream_readdata),
      .SS_OCT_SOPC_burst_0_upstream_readdata_from_sa                                             (SS_OCT_SOPC_burst_0_upstream_readdata_from_sa),
      .SS_OCT_SOPC_burst_0_upstream_readdatavalid                                                (SS_OCT_SOPC_burst_0_upstream_readdatavalid),
      .SS_OCT_SOPC_burst_0_upstream_waitrequest                                                  (SS_OCT_SOPC_burst_0_upstream_waitrequest),
      .SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa                                          (SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa),
      .SS_OCT_SOPC_burst_0_upstream_write                                                        (SS_OCT_SOPC_burst_0_upstream_write),
      .SS_OCT_SOPC_burst_0_upstream_writedata                                                    (SS_OCT_SOPC_burst_0_upstream_writedata),
      .clk                                                                                       (ddr2_phy_clk_out),
      .clock_crossing_master_ddr2_m1_address_to_slave                                            (clock_crossing_master_ddr2_m1_address_to_slave),
      .clock_crossing_master_ddr2_m1_burstcount                                                  (clock_crossing_master_ddr2_m1_burstcount),
      .clock_crossing_master_ddr2_m1_byteenable                                                  (clock_crossing_master_ddr2_m1_byteenable),
      .clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream                        (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_latency_counter                                             (clock_crossing_master_ddr2_m1_latency_counter),
      .clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream              (clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_read                                                        (clock_crossing_master_ddr2_m1_read),
      .clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream                (clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register (clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register),
      .clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream                       (clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_write                                                       (clock_crossing_master_ddr2_m1_write),
      .clock_crossing_master_ddr2_m1_writedata                                                   (clock_crossing_master_ddr2_m1_writedata),
      .d1_SS_OCT_SOPC_burst_0_upstream_end_xfer                                                  (d1_SS_OCT_SOPC_burst_0_upstream_end_xfer),
      .reset_n                                                                                   (ddr2_phy_clk_out_reset_n)
    );

  SS_OCT_SOPC_burst_0_downstream_arbitrator the_SS_OCT_SOPC_burst_0_downstream
    (
      .SS_OCT_SOPC_burst_0_downstream_address                                (SS_OCT_SOPC_burst_0_downstream_address),
      .SS_OCT_SOPC_burst_0_downstream_address_to_slave                       (SS_OCT_SOPC_burst_0_downstream_address_to_slave),
      .SS_OCT_SOPC_burst_0_downstream_burstcount                             (SS_OCT_SOPC_burst_0_downstream_burstcount),
      .SS_OCT_SOPC_burst_0_downstream_byteenable                             (SS_OCT_SOPC_burst_0_downstream_byteenable),
      .SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1                        (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_latency_counter                        (SS_OCT_SOPC_burst_0_downstream_latency_counter),
      .SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1              (SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_read                                   (SS_OCT_SOPC_burst_0_downstream_read),
      .SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1                (SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register (SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register),
      .SS_OCT_SOPC_burst_0_downstream_readdata                               (SS_OCT_SOPC_burst_0_downstream_readdata),
      .SS_OCT_SOPC_burst_0_downstream_readdatavalid                          (SS_OCT_SOPC_burst_0_downstream_readdatavalid),
      .SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1                       (SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_reset_n                                (SS_OCT_SOPC_burst_0_downstream_reset_n),
      .SS_OCT_SOPC_burst_0_downstream_waitrequest                            (SS_OCT_SOPC_burst_0_downstream_waitrequest),
      .SS_OCT_SOPC_burst_0_downstream_write                                  (SS_OCT_SOPC_burst_0_downstream_write),
      .SS_OCT_SOPC_burst_0_downstream_writedata                              (SS_OCT_SOPC_burst_0_downstream_writedata),
      .clk                                                                   (ddr2_phy_clk_out),
      .d1_ddr2_s1_end_xfer                                                   (d1_ddr2_s1_end_xfer),
      .ddr2_s1_readdata_from_sa                                              (ddr2_s1_readdata_from_sa),
      .ddr2_s1_waitrequest_n_from_sa                                         (ddr2_s1_waitrequest_n_from_sa),
      .reset_n                                                               (ddr2_phy_clk_out_reset_n)
    );

  SS_OCT_SOPC_burst_0 the_SS_OCT_SOPC_burst_0
    (
      .clk                         (ddr2_phy_clk_out),
      .downstream_address          (SS_OCT_SOPC_burst_0_downstream_address),
      .downstream_arbitrationshare (SS_OCT_SOPC_burst_0_downstream_arbitrationshare),
      .downstream_burstcount       (SS_OCT_SOPC_burst_0_downstream_burstcount),
      .downstream_byteenable       (SS_OCT_SOPC_burst_0_downstream_byteenable),
      .downstream_debugaccess      (SS_OCT_SOPC_burst_0_downstream_debugaccess),
      .downstream_nativeaddress    (SS_OCT_SOPC_burst_0_downstream_nativeaddress),
      .downstream_read             (SS_OCT_SOPC_burst_0_downstream_read),
      .downstream_readdata         (SS_OCT_SOPC_burst_0_downstream_readdata),
      .downstream_readdatavalid    (SS_OCT_SOPC_burst_0_downstream_readdatavalid),
      .downstream_waitrequest      (SS_OCT_SOPC_burst_0_downstream_waitrequest),
      .downstream_write            (SS_OCT_SOPC_burst_0_downstream_write),
      .downstream_writedata        (SS_OCT_SOPC_burst_0_downstream_writedata),
      .reset_n                     (SS_OCT_SOPC_burst_0_downstream_reset_n),
      .upstream_address            (SS_OCT_SOPC_burst_0_upstream_byteaddress),
      .upstream_burstcount         (SS_OCT_SOPC_burst_0_upstream_burstcount),
      .upstream_byteenable         (SS_OCT_SOPC_burst_0_upstream_byteenable),
      .upstream_debugaccess        (SS_OCT_SOPC_burst_0_upstream_debugaccess),
      .upstream_nativeaddress      (SS_OCT_SOPC_burst_0_upstream_address),
      .upstream_read               (SS_OCT_SOPC_burst_0_upstream_read),
      .upstream_readdata           (SS_OCT_SOPC_burst_0_upstream_readdata),
      .upstream_readdatavalid      (SS_OCT_SOPC_burst_0_upstream_readdatavalid),
      .upstream_waitrequest        (SS_OCT_SOPC_burst_0_upstream_waitrequest),
      .upstream_write              (SS_OCT_SOPC_burst_0_upstream_write),
      .upstream_writedata          (SS_OCT_SOPC_burst_0_upstream_writedata)
    );

  SS_OCT_SOPC_clock_0_in_arbitrator the_SS_OCT_SOPC_clock_0_in
    (
      .SS_OCT_SOPC_clock_0_in_address                                            (SS_OCT_SOPC_clock_0_in_address),
      .SS_OCT_SOPC_clock_0_in_byteenable                                         (SS_OCT_SOPC_clock_0_in_byteenable),
      .SS_OCT_SOPC_clock_0_in_endofpacket                                        (SS_OCT_SOPC_clock_0_in_endofpacket),
      .SS_OCT_SOPC_clock_0_in_endofpacket_from_sa                                (SS_OCT_SOPC_clock_0_in_endofpacket_from_sa),
      .SS_OCT_SOPC_clock_0_in_nativeaddress                                      (SS_OCT_SOPC_clock_0_in_nativeaddress),
      .SS_OCT_SOPC_clock_0_in_read                                               (SS_OCT_SOPC_clock_0_in_read),
      .SS_OCT_SOPC_clock_0_in_readdata                                           (SS_OCT_SOPC_clock_0_in_readdata),
      .SS_OCT_SOPC_clock_0_in_readdata_from_sa                                   (SS_OCT_SOPC_clock_0_in_readdata_from_sa),
      .SS_OCT_SOPC_clock_0_in_reset_n                                            (SS_OCT_SOPC_clock_0_in_reset_n),
      .SS_OCT_SOPC_clock_0_in_waitrequest                                        (SS_OCT_SOPC_clock_0_in_waitrequest),
      .SS_OCT_SOPC_clock_0_in_waitrequest_from_sa                                (SS_OCT_SOPC_clock_0_in_waitrequest_from_sa),
      .SS_OCT_SOPC_clock_0_in_write                                              (SS_OCT_SOPC_clock_0_in_write),
      .SS_OCT_SOPC_clock_0_in_writedata                                          (SS_OCT_SOPC_clock_0_in_writedata),
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_granted_SS_OCT_SOPC_clock_0_in                            (cpu_data_master_granted_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in                  (cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in                    (cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_requests_SS_OCT_SOPC_clock_0_in                           (cpu_data_master_requests_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_SS_OCT_SOPC_clock_0_in_end_xfer                                        (d1_SS_OCT_SOPC_clock_0_in_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  SS_OCT_SOPC_clock_0_out_arbitrator the_SS_OCT_SOPC_clock_0_out
    (
      .SS_OCT_SOPC_clock_0_out_address                  (SS_OCT_SOPC_clock_0_out_address),
      .SS_OCT_SOPC_clock_0_out_address_to_slave         (SS_OCT_SOPC_clock_0_out_address_to_slave),
      .SS_OCT_SOPC_clock_0_out_byteenable               (SS_OCT_SOPC_clock_0_out_byteenable),
      .SS_OCT_SOPC_clock_0_out_granted_pll_s1           (SS_OCT_SOPC_clock_0_out_granted_pll_s1),
      .SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1 (SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1),
      .SS_OCT_SOPC_clock_0_out_read                     (SS_OCT_SOPC_clock_0_out_read),
      .SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1   (SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1),
      .SS_OCT_SOPC_clock_0_out_readdata                 (SS_OCT_SOPC_clock_0_out_readdata),
      .SS_OCT_SOPC_clock_0_out_requests_pll_s1          (SS_OCT_SOPC_clock_0_out_requests_pll_s1),
      .SS_OCT_SOPC_clock_0_out_reset_n                  (SS_OCT_SOPC_clock_0_out_reset_n),
      .SS_OCT_SOPC_clock_0_out_waitrequest              (SS_OCT_SOPC_clock_0_out_waitrequest),
      .SS_OCT_SOPC_clock_0_out_write                    (SS_OCT_SOPC_clock_0_out_write),
      .SS_OCT_SOPC_clock_0_out_writedata                (SS_OCT_SOPC_clock_0_out_writedata),
      .clk                                              (clk_50),
      .d1_pll_s1_end_xfer                               (d1_pll_s1_end_xfer),
      .pll_s1_readdata_from_sa                          (pll_s1_readdata_from_sa),
      .reset_n                                          (clk_50_reset_n)
    );

  SS_OCT_SOPC_clock_0 the_SS_OCT_SOPC_clock_0
    (
      .master_address       (SS_OCT_SOPC_clock_0_out_address),
      .master_byteenable    (SS_OCT_SOPC_clock_0_out_byteenable),
      .master_clk           (clk_50),
      .master_endofpacket   (SS_OCT_SOPC_clock_0_out_endofpacket),
      .master_nativeaddress (SS_OCT_SOPC_clock_0_out_nativeaddress),
      .master_read          (SS_OCT_SOPC_clock_0_out_read),
      .master_readdata      (SS_OCT_SOPC_clock_0_out_readdata),
      .master_reset_n       (SS_OCT_SOPC_clock_0_out_reset_n),
      .master_waitrequest   (SS_OCT_SOPC_clock_0_out_waitrequest),
      .master_write         (SS_OCT_SOPC_clock_0_out_write),
      .master_writedata     (SS_OCT_SOPC_clock_0_out_writedata),
      .slave_address        (SS_OCT_SOPC_clock_0_in_address),
      .slave_byteenable     (SS_OCT_SOPC_clock_0_in_byteenable),
      .slave_clk            (pll_sys_clk),
      .slave_endofpacket    (SS_OCT_SOPC_clock_0_in_endofpacket),
      .slave_nativeaddress  (SS_OCT_SOPC_clock_0_in_nativeaddress),
      .slave_read           (SS_OCT_SOPC_clock_0_in_read),
      .slave_readdata       (SS_OCT_SOPC_clock_0_in_readdata),
      .slave_reset_n        (SS_OCT_SOPC_clock_0_in_reset_n),
      .slave_waitrequest    (SS_OCT_SOPC_clock_0_in_waitrequest),
      .slave_write          (SS_OCT_SOPC_clock_0_in_write),
      .slave_writedata      (SS_OCT_SOPC_clock_0_in_writedata)
    );

  clock_crossing_ddr2_cpu_s1_arbitrator the_clock_crossing_ddr2_cpu_s1
    (
      .clk                                                                       (pll_sys_clk),
      .clock_crossing_ddr2_cpu_s1_address                                        (clock_crossing_ddr2_cpu_s1_address),
      .clock_crossing_ddr2_cpu_s1_byteenable                                     (clock_crossing_ddr2_cpu_s1_byteenable),
      .clock_crossing_ddr2_cpu_s1_endofpacket                                    (clock_crossing_ddr2_cpu_s1_endofpacket),
      .clock_crossing_ddr2_cpu_s1_endofpacket_from_sa                            (clock_crossing_ddr2_cpu_s1_endofpacket_from_sa),
      .clock_crossing_ddr2_cpu_s1_nativeaddress                                  (clock_crossing_ddr2_cpu_s1_nativeaddress),
      .clock_crossing_ddr2_cpu_s1_read                                           (clock_crossing_ddr2_cpu_s1_read),
      .clock_crossing_ddr2_cpu_s1_readdata                                       (clock_crossing_ddr2_cpu_s1_readdata),
      .clock_crossing_ddr2_cpu_s1_readdata_from_sa                               (clock_crossing_ddr2_cpu_s1_readdata_from_sa),
      .clock_crossing_ddr2_cpu_s1_readdatavalid                                  (clock_crossing_ddr2_cpu_s1_readdatavalid),
      .clock_crossing_ddr2_cpu_s1_reset_n                                        (clock_crossing_ddr2_cpu_s1_reset_n),
      .clock_crossing_ddr2_cpu_s1_waitrequest                                    (clock_crossing_ddr2_cpu_s1_waitrequest),
      .clock_crossing_ddr2_cpu_s1_waitrequest_from_sa                            (clock_crossing_ddr2_cpu_s1_waitrequest_from_sa),
      .clock_crossing_ddr2_cpu_s1_write                                          (clock_crossing_ddr2_cpu_s1_write),
      .clock_crossing_ddr2_cpu_s1_writedata                                      (clock_crossing_ddr2_cpu_s1_writedata),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_granted_clock_crossing_ddr2_cpu_s1                        (cpu_data_master_granted_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1              (cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1                (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_requests_clock_crossing_ddr2_cpu_s1                       (cpu_data_master_requests_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_clock_crossing_ddr2_cpu_s1_end_xfer                                    (d1_clock_crossing_ddr2_cpu_s1_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  clock_crossing_ddr2_cpu_m1_arbitrator the_clock_crossing_ddr2_cpu_m1
    (
      .clk                                                                               (ddr2_phy_clk_out),
      .clock_crossing_ddr2_cpu_m1_address                                                (clock_crossing_ddr2_cpu_m1_address),
      .clock_crossing_ddr2_cpu_m1_address_to_slave                                       (clock_crossing_ddr2_cpu_m1_address_to_slave),
      .clock_crossing_ddr2_cpu_m1_byteenable                                             (clock_crossing_ddr2_cpu_m1_byteenable),
      .clock_crossing_ddr2_cpu_m1_endofpacket                                            (clock_crossing_ddr2_cpu_m1_endofpacket),
      .clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1                        (clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_latency_counter                                        (clock_crossing_ddr2_cpu_m1_latency_counter),
      .clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1              (clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_read                                                   (clock_crossing_ddr2_cpu_m1_read),
      .clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1                (clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register (clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register),
      .clock_crossing_ddr2_cpu_m1_readdata                                               (clock_crossing_ddr2_cpu_m1_readdata),
      .clock_crossing_ddr2_cpu_m1_readdatavalid                                          (clock_crossing_ddr2_cpu_m1_readdatavalid),
      .clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1                       (clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_reset_n                                                (clock_crossing_ddr2_cpu_m1_reset_n),
      .clock_crossing_ddr2_cpu_m1_waitrequest                                            (clock_crossing_ddr2_cpu_m1_waitrequest),
      .clock_crossing_ddr2_cpu_m1_write                                                  (clock_crossing_ddr2_cpu_m1_write),
      .clock_crossing_ddr2_cpu_m1_writedata                                              (clock_crossing_ddr2_cpu_m1_writedata),
      .d1_pipeline_bridge_ddr2_s1_end_xfer                                               (d1_pipeline_bridge_ddr2_s1_end_xfer),
      .pipeline_bridge_ddr2_s1_endofpacket_from_sa                                       (pipeline_bridge_ddr2_s1_endofpacket_from_sa),
      .pipeline_bridge_ddr2_s1_readdata_from_sa                                          (pipeline_bridge_ddr2_s1_readdata_from_sa),
      .pipeline_bridge_ddr2_s1_waitrequest_from_sa                                       (pipeline_bridge_ddr2_s1_waitrequest_from_sa),
      .reset_n                                                                           (ddr2_phy_clk_out_reset_n)
    );

  clock_crossing_ddr2_cpu the_clock_crossing_ddr2_cpu
    (
      .master_address       (clock_crossing_ddr2_cpu_m1_address),
      .master_byteenable    (clock_crossing_ddr2_cpu_m1_byteenable),
      .master_clk           (ddr2_phy_clk_out),
      .master_endofpacket   (clock_crossing_ddr2_cpu_m1_endofpacket),
      .master_nativeaddress (clock_crossing_ddr2_cpu_m1_nativeaddress),
      .master_read          (clock_crossing_ddr2_cpu_m1_read),
      .master_readdata      (clock_crossing_ddr2_cpu_m1_readdata),
      .master_readdatavalid (clock_crossing_ddr2_cpu_m1_readdatavalid),
      .master_reset_n       (clock_crossing_ddr2_cpu_m1_reset_n),
      .master_waitrequest   (clock_crossing_ddr2_cpu_m1_waitrequest),
      .master_write         (clock_crossing_ddr2_cpu_m1_write),
      .master_writedata     (clock_crossing_ddr2_cpu_m1_writedata),
      .slave_address        (clock_crossing_ddr2_cpu_s1_address),
      .slave_byteenable     (clock_crossing_ddr2_cpu_s1_byteenable),
      .slave_clk            (pll_sys_clk),
      .slave_endofpacket    (clock_crossing_ddr2_cpu_s1_endofpacket),
      .slave_nativeaddress  (clock_crossing_ddr2_cpu_s1_nativeaddress),
      .slave_read           (clock_crossing_ddr2_cpu_s1_read),
      .slave_readdata       (clock_crossing_ddr2_cpu_s1_readdata),
      .slave_readdatavalid  (clock_crossing_ddr2_cpu_s1_readdatavalid),
      .slave_reset_n        (clock_crossing_ddr2_cpu_s1_reset_n),
      .slave_waitrequest    (clock_crossing_ddr2_cpu_s1_waitrequest),
      .slave_write          (clock_crossing_ddr2_cpu_s1_write),
      .slave_writedata      (clock_crossing_ddr2_cpu_s1_writedata)
    );

  clock_crossing_master_ddr2_s1_arbitrator the_clock_crossing_master_ddr2_s1
    (
      .clk                                                                      (clk_50),
      .clock_crossing_master_ddr2_s1_address                                    (clock_crossing_master_ddr2_s1_address),
      .clock_crossing_master_ddr2_s1_burstcount                                 (clock_crossing_master_ddr2_s1_burstcount),
      .clock_crossing_master_ddr2_s1_byteenable                                 (clock_crossing_master_ddr2_s1_byteenable),
      .clock_crossing_master_ddr2_s1_endofpacket                                (clock_crossing_master_ddr2_s1_endofpacket),
      .clock_crossing_master_ddr2_s1_endofpacket_from_sa                        (clock_crossing_master_ddr2_s1_endofpacket_from_sa),
      .clock_crossing_master_ddr2_s1_nativeaddress                              (clock_crossing_master_ddr2_s1_nativeaddress),
      .clock_crossing_master_ddr2_s1_read                                       (clock_crossing_master_ddr2_s1_read),
      .clock_crossing_master_ddr2_s1_readdata                                   (clock_crossing_master_ddr2_s1_readdata),
      .clock_crossing_master_ddr2_s1_readdata_from_sa                           (clock_crossing_master_ddr2_s1_readdata_from_sa),
      .clock_crossing_master_ddr2_s1_readdatavalid                              (clock_crossing_master_ddr2_s1_readdatavalid),
      .clock_crossing_master_ddr2_s1_reset_n                                    (clock_crossing_master_ddr2_s1_reset_n),
      .clock_crossing_master_ddr2_s1_waitrequest                                (clock_crossing_master_ddr2_s1_waitrequest),
      .clock_crossing_master_ddr2_s1_waitrequest_from_sa                        (clock_crossing_master_ddr2_s1_waitrequest_from_sa),
      .clock_crossing_master_ddr2_s1_write                                      (clock_crossing_master_ddr2_s1_write),
      .clock_crossing_master_ddr2_s1_writedata                                  (clock_crossing_master_ddr2_s1_writedata),
      .d1_clock_crossing_master_ddr2_s1_end_xfer                                (d1_clock_crossing_master_ddr2_s1_end_xfer),
      .master_read_avalon_master_address_to_slave                               (master_read_avalon_master_address_to_slave),
      .master_read_avalon_master_burstcount                                     (master_read_avalon_master_burstcount),
      .master_read_avalon_master_read                                           (master_read_avalon_master_read),
      .master_read_granted_clock_crossing_master_ddr2_s1                        (master_read_granted_clock_crossing_master_ddr2_s1),
      .master_read_latency_counter                                              (master_read_latency_counter),
      .master_read_qualified_request_clock_crossing_master_ddr2_s1              (master_read_qualified_request_clock_crossing_master_ddr2_s1),
      .master_read_read_data_valid_clock_crossing_master_ddr2_s1                (master_read_read_data_valid_clock_crossing_master_ddr2_s1),
      .master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register (master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register),
      .master_read_requests_clock_crossing_master_ddr2_s1                       (master_read_requests_clock_crossing_master_ddr2_s1),
      .master_write_avalon_master_address_to_slave                              (master_write_avalon_master_address_to_slave),
      .master_write_avalon_master_burstcount                                    (master_write_avalon_master_burstcount),
      .master_write_avalon_master_byteenable                                    (master_write_avalon_master_byteenable),
      .master_write_avalon_master_write                                         (master_write_avalon_master_write),
      .master_write_avalon_master_writedata                                     (master_write_avalon_master_writedata),
      .master_write_granted_clock_crossing_master_ddr2_s1                       (master_write_granted_clock_crossing_master_ddr2_s1),
      .master_write_qualified_request_clock_crossing_master_ddr2_s1             (master_write_qualified_request_clock_crossing_master_ddr2_s1),
      .master_write_requests_clock_crossing_master_ddr2_s1                      (master_write_requests_clock_crossing_master_ddr2_s1),
      .reset_n                                                                  (clk_50_reset_n)
    );

  clock_crossing_master_ddr2_m1_arbitrator the_clock_crossing_master_ddr2_m1
    (
      .SS_OCT_SOPC_burst_0_upstream_readdata_from_sa                                             (SS_OCT_SOPC_burst_0_upstream_readdata_from_sa),
      .SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa                                          (SS_OCT_SOPC_burst_0_upstream_waitrequest_from_sa),
      .clk                                                                                       (ddr2_phy_clk_out),
      .clock_crossing_master_ddr2_m1_address                                                     (clock_crossing_master_ddr2_m1_address),
      .clock_crossing_master_ddr2_m1_address_to_slave                                            (clock_crossing_master_ddr2_m1_address_to_slave),
      .clock_crossing_master_ddr2_m1_burstcount                                                  (clock_crossing_master_ddr2_m1_burstcount),
      .clock_crossing_master_ddr2_m1_byteenable                                                  (clock_crossing_master_ddr2_m1_byteenable),
      .clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream                        (clock_crossing_master_ddr2_m1_granted_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_latency_counter                                             (clock_crossing_master_ddr2_m1_latency_counter),
      .clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream              (clock_crossing_master_ddr2_m1_qualified_request_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_read                                                        (clock_crossing_master_ddr2_m1_read),
      .clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream                (clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register (clock_crossing_master_ddr2_m1_read_data_valid_SS_OCT_SOPC_burst_0_upstream_shift_register),
      .clock_crossing_master_ddr2_m1_readdata                                                    (clock_crossing_master_ddr2_m1_readdata),
      .clock_crossing_master_ddr2_m1_readdatavalid                                               (clock_crossing_master_ddr2_m1_readdatavalid),
      .clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream                       (clock_crossing_master_ddr2_m1_requests_SS_OCT_SOPC_burst_0_upstream),
      .clock_crossing_master_ddr2_m1_reset_n                                                     (clock_crossing_master_ddr2_m1_reset_n),
      .clock_crossing_master_ddr2_m1_waitrequest                                                 (clock_crossing_master_ddr2_m1_waitrequest),
      .clock_crossing_master_ddr2_m1_write                                                       (clock_crossing_master_ddr2_m1_write),
      .clock_crossing_master_ddr2_m1_writedata                                                   (clock_crossing_master_ddr2_m1_writedata),
      .d1_SS_OCT_SOPC_burst_0_upstream_end_xfer                                                  (d1_SS_OCT_SOPC_burst_0_upstream_end_xfer),
      .reset_n                                                                                   (ddr2_phy_clk_out_reset_n)
    );

  clock_crossing_master_ddr2 the_clock_crossing_master_ddr2
    (
      .master_address       (clock_crossing_master_ddr2_m1_address),
      .master_burstcount    (clock_crossing_master_ddr2_m1_burstcount),
      .master_byteenable    (clock_crossing_master_ddr2_m1_byteenable),
      .master_clk           (ddr2_phy_clk_out),
      .master_endofpacket   (clock_crossing_master_ddr2_m1_endofpacket),
      .master_nativeaddress (clock_crossing_master_ddr2_m1_nativeaddress),
      .master_read          (clock_crossing_master_ddr2_m1_read),
      .master_readdata      (clock_crossing_master_ddr2_m1_readdata),
      .master_readdatavalid (clock_crossing_master_ddr2_m1_readdatavalid),
      .master_reset_n       (clock_crossing_master_ddr2_m1_reset_n),
      .master_waitrequest   (clock_crossing_master_ddr2_m1_waitrequest),
      .master_write         (clock_crossing_master_ddr2_m1_write),
      .master_writedata     (clock_crossing_master_ddr2_m1_writedata),
      .slave_address        (clock_crossing_master_ddr2_s1_address),
      .slave_burstcount     (clock_crossing_master_ddr2_s1_burstcount),
      .slave_byteenable     (clock_crossing_master_ddr2_s1_byteenable),
      .slave_clk            (clk_50),
      .slave_endofpacket    (clock_crossing_master_ddr2_s1_endofpacket),
      .slave_nativeaddress  (clock_crossing_master_ddr2_s1_nativeaddress),
      .slave_read           (clock_crossing_master_ddr2_s1_read),
      .slave_readdata       (clock_crossing_master_ddr2_s1_readdata),
      .slave_readdatavalid  (clock_crossing_master_ddr2_s1_readdatavalid),
      .slave_reset_n        (clock_crossing_master_ddr2_s1_reset_n),
      .slave_waitrequest    (clock_crossing_master_ddr2_s1_waitrequest),
      .slave_write          (clock_crossing_master_ddr2_s1_write),
      .slave_writedata      (clock_crossing_master_ddr2_s1_writedata)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                               (cpu_data_master_debugaccess),
      .cpu_data_master_granted_cpu_jtag_debug_module                             (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module                   (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                     (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_requests_cpu_jtag_debug_module                            (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                   (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_jtag_debug_module                      (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_latency_counter                                    (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module            (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_read                                               (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module              (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_requests_cpu_jtag_debug_module                     (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_jtag_debug_module_address                                             (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                                       (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                                          (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                                          (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                                         (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                            (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                                    (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                                             (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                                        (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                                (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                               (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                           (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                                         (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .SS_OCT_SOPC_clock_0_in_readdata_from_sa                                   (SS_OCT_SOPC_clock_0_in_readdata_from_sa),
      .SS_OCT_SOPC_clock_0_in_waitrequest_from_sa                                (SS_OCT_SOPC_clock_0_in_waitrequest_from_sa),
      .clk                                                                       (pll_sys_clk),
      .clock_crossing_ddr2_cpu_s1_readdata_from_sa                               (clock_crossing_ddr2_cpu_s1_readdata_from_sa),
      .clock_crossing_ddr2_cpu_s1_waitrequest_from_sa                            (clock_crossing_ddr2_cpu_s1_waitrequest_from_sa),
      .cpu_data_master_address                                                   (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_byteenable_ext_flash_s1                                   (cpu_data_master_byteenable_ext_flash_s1),
      .cpu_data_master_dbs_address                                               (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_16                                              (cpu_data_master_dbs_write_16),
      .cpu_data_master_granted_SS_OCT_SOPC_clock_0_in                            (cpu_data_master_granted_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_granted_clock_crossing_ddr2_cpu_s1                        (cpu_data_master_granted_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_granted_cpu_jtag_debug_module                             (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_granted_descriptor_memory_s1                              (cpu_data_master_granted_descriptor_memory_s1),
      .cpu_data_master_granted_ext_flash_s1                                      (cpu_data_master_granted_ext_flash_s1),
      .cpu_data_master_granted_high_res_timer_s1                                 (cpu_data_master_granted_high_res_timer_s1),
      .cpu_data_master_granted_jtag_uart_avalon_jtag_slave                       (cpu_data_master_granted_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_granted_onchip_memory_s1                                  (cpu_data_master_granted_onchip_memory_s1),
      .cpu_data_master_granted_packet_memory_s1                                  (cpu_data_master_granted_packet_memory_s1),
      .cpu_data_master_granted_sgdma_rx_csr                                      (cpu_data_master_granted_sgdma_rx_csr),
      .cpu_data_master_granted_sgdma_tx_csr                                      (cpu_data_master_granted_sgdma_tx_csr),
      .cpu_data_master_granted_sys_timer_s1                                      (cpu_data_master_granted_sys_timer_s1),
      .cpu_data_master_granted_sysid_control_slave                               (cpu_data_master_granted_sysid_control_slave),
      .cpu_data_master_granted_tse_mac_control_port                              (cpu_data_master_granted_tse_mac_control_port),
      .cpu_data_master_granted_vol_recording_done_pio_s1                         (cpu_data_master_granted_vol_recording_done_pio_s1),
      .cpu_data_master_granted_vol_transfer_done_pio_s1                          (cpu_data_master_granted_vol_transfer_done_pio_s1),
      .cpu_data_master_irq                                                       (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in                  (cpu_data_master_qualified_request_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1              (cpu_data_master_qualified_request_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module                   (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_qualified_request_descriptor_memory_s1                    (cpu_data_master_qualified_request_descriptor_memory_s1),
      .cpu_data_master_qualified_request_ext_flash_s1                            (cpu_data_master_qualified_request_ext_flash_s1),
      .cpu_data_master_qualified_request_high_res_timer_s1                       (cpu_data_master_qualified_request_high_res_timer_s1),
      .cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave             (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_qualified_request_onchip_memory_s1                        (cpu_data_master_qualified_request_onchip_memory_s1),
      .cpu_data_master_qualified_request_packet_memory_s1                        (cpu_data_master_qualified_request_packet_memory_s1),
      .cpu_data_master_qualified_request_sgdma_rx_csr                            (cpu_data_master_qualified_request_sgdma_rx_csr),
      .cpu_data_master_qualified_request_sgdma_tx_csr                            (cpu_data_master_qualified_request_sgdma_tx_csr),
      .cpu_data_master_qualified_request_sys_timer_s1                            (cpu_data_master_qualified_request_sys_timer_s1),
      .cpu_data_master_qualified_request_sysid_control_slave                     (cpu_data_master_qualified_request_sysid_control_slave),
      .cpu_data_master_qualified_request_tse_mac_control_port                    (cpu_data_master_qualified_request_tse_mac_control_port),
      .cpu_data_master_qualified_request_vol_recording_done_pio_s1               (cpu_data_master_qualified_request_vol_recording_done_pio_s1),
      .cpu_data_master_qualified_request_vol_transfer_done_pio_s1                (cpu_data_master_qualified_request_vol_transfer_done_pio_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in                    (cpu_data_master_read_data_valid_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1                (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                     (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_descriptor_memory_s1                      (cpu_data_master_read_data_valid_descriptor_memory_s1),
      .cpu_data_master_read_data_valid_ext_flash_s1                              (cpu_data_master_read_data_valid_ext_flash_s1),
      .cpu_data_master_read_data_valid_high_res_timer_s1                         (cpu_data_master_read_data_valid_high_res_timer_s1),
      .cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave               (cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_read_data_valid_onchip_memory_s1                          (cpu_data_master_read_data_valid_onchip_memory_s1),
      .cpu_data_master_read_data_valid_packet_memory_s1                          (cpu_data_master_read_data_valid_packet_memory_s1),
      .cpu_data_master_read_data_valid_sgdma_rx_csr                              (cpu_data_master_read_data_valid_sgdma_rx_csr),
      .cpu_data_master_read_data_valid_sgdma_tx_csr                              (cpu_data_master_read_data_valid_sgdma_tx_csr),
      .cpu_data_master_read_data_valid_sys_timer_s1                              (cpu_data_master_read_data_valid_sys_timer_s1),
      .cpu_data_master_read_data_valid_sysid_control_slave                       (cpu_data_master_read_data_valid_sysid_control_slave),
      .cpu_data_master_read_data_valid_tse_mac_control_port                      (cpu_data_master_read_data_valid_tse_mac_control_port),
      .cpu_data_master_read_data_valid_vol_recording_done_pio_s1                 (cpu_data_master_read_data_valid_vol_recording_done_pio_s1),
      .cpu_data_master_read_data_valid_vol_transfer_done_pio_s1                  (cpu_data_master_read_data_valid_vol_transfer_done_pio_s1),
      .cpu_data_master_readdata                                                  (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                             (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_SS_OCT_SOPC_clock_0_in                           (cpu_data_master_requests_SS_OCT_SOPC_clock_0_in),
      .cpu_data_master_requests_clock_crossing_ddr2_cpu_s1                       (cpu_data_master_requests_clock_crossing_ddr2_cpu_s1),
      .cpu_data_master_requests_cpu_jtag_debug_module                            (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_requests_descriptor_memory_s1                             (cpu_data_master_requests_descriptor_memory_s1),
      .cpu_data_master_requests_ext_flash_s1                                     (cpu_data_master_requests_ext_flash_s1),
      .cpu_data_master_requests_high_res_timer_s1                                (cpu_data_master_requests_high_res_timer_s1),
      .cpu_data_master_requests_jtag_uart_avalon_jtag_slave                      (cpu_data_master_requests_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_requests_onchip_memory_s1                                 (cpu_data_master_requests_onchip_memory_s1),
      .cpu_data_master_requests_packet_memory_s1                                 (cpu_data_master_requests_packet_memory_s1),
      .cpu_data_master_requests_sgdma_rx_csr                                     (cpu_data_master_requests_sgdma_rx_csr),
      .cpu_data_master_requests_sgdma_tx_csr                                     (cpu_data_master_requests_sgdma_tx_csr),
      .cpu_data_master_requests_sys_timer_s1                                     (cpu_data_master_requests_sys_timer_s1),
      .cpu_data_master_requests_sysid_control_slave                              (cpu_data_master_requests_sysid_control_slave),
      .cpu_data_master_requests_tse_mac_control_port                             (cpu_data_master_requests_tse_mac_control_port),
      .cpu_data_master_requests_vol_recording_done_pio_s1                        (cpu_data_master_requests_vol_recording_done_pio_s1),
      .cpu_data_master_requests_vol_transfer_done_pio_s1                         (cpu_data_master_requests_vol_transfer_done_pio_s1),
      .cpu_data_master_waitrequest                                               (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .cpu_jtag_debug_module_readdata_from_sa                                    (cpu_jtag_debug_module_readdata_from_sa),
      .d1_SS_OCT_SOPC_clock_0_in_end_xfer                                        (d1_SS_OCT_SOPC_clock_0_in_end_xfer),
      .d1_clock_crossing_ddr2_cpu_s1_end_xfer                                    (d1_clock_crossing_ddr2_cpu_s1_end_xfer),
      .d1_cpu_jtag_debug_module_end_xfer                                         (d1_cpu_jtag_debug_module_end_xfer),
      .d1_descriptor_memory_s1_end_xfer                                          (d1_descriptor_memory_s1_end_xfer),
      .d1_flash_tristate_bridge_avalon_slave_end_xfer                            (d1_flash_tristate_bridge_avalon_slave_end_xfer),
      .d1_high_res_timer_s1_end_xfer                                             (d1_high_res_timer_s1_end_xfer),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                   (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_onchip_memory_s1_end_xfer                                              (d1_onchip_memory_s1_end_xfer),
      .d1_packet_memory_s1_end_xfer                                              (d1_packet_memory_s1_end_xfer),
      .d1_sgdma_rx_csr_end_xfer                                                  (d1_sgdma_rx_csr_end_xfer),
      .d1_sgdma_tx_csr_end_xfer                                                  (d1_sgdma_tx_csr_end_xfer),
      .d1_sys_timer_s1_end_xfer                                                  (d1_sys_timer_s1_end_xfer),
      .d1_sysid_control_slave_end_xfer                                           (d1_sysid_control_slave_end_xfer),
      .d1_tse_mac_control_port_end_xfer                                          (d1_tse_mac_control_port_end_xfer),
      .d1_vol_recording_done_pio_s1_end_xfer                                     (d1_vol_recording_done_pio_s1_end_xfer),
      .d1_vol_transfer_done_pio_s1_end_xfer                                      (d1_vol_transfer_done_pio_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                                     (descriptor_memory_s1_readdata_from_sa),
      .ext_flash_s1_wait_counter_eq_0                                            (ext_flash_s1_wait_counter_eq_0),
      .high_res_timer_s1_irq_from_sa                                             (high_res_timer_s1_irq_from_sa),
      .high_res_timer_s1_readdata_from_sa                                        (high_res_timer_s1_readdata_from_sa),
      .incoming_flash_tristate_bridge_data_with_Xs_converted_to_0                (incoming_flash_tristate_bridge_data_with_Xs_converted_to_0),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                   (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                              (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                           (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .onchip_memory_s1_readdata_from_sa                                         (onchip_memory_s1_readdata_from_sa),
      .packet_memory_s1_readdata_from_sa                                         (packet_memory_s1_readdata_from_sa),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sgdma_rx_csr_irq_from_sa                                                  (sgdma_rx_csr_irq_from_sa),
      .sgdma_rx_csr_readdata_from_sa                                             (sgdma_rx_csr_readdata_from_sa),
      .sgdma_tx_csr_irq_from_sa                                                  (sgdma_tx_csr_irq_from_sa),
      .sgdma_tx_csr_readdata_from_sa                                             (sgdma_tx_csr_readdata_from_sa),
      .sys_timer_s1_irq_from_sa                                                  (sys_timer_s1_irq_from_sa),
      .sys_timer_s1_readdata_from_sa                                             (sys_timer_s1_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                      (sysid_control_slave_readdata_from_sa),
      .tse_mac_control_port_readdata_from_sa                                     (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_waitrequest_from_sa                                  (tse_mac_control_port_waitrequest_from_sa),
      .vol_recording_done_pio_s1_readdata_from_sa                                (vol_recording_done_pio_s1_readdata_from_sa),
      .vol_transfer_done_pio_s1_readdata_from_sa                                 (vol_transfer_done_pio_s1_readdata_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                            (pll_sys_clk),
      .cpu_instruction_master_address                                 (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                        (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_dbs_address                             (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_cpu_jtag_debug_module           (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_granted_descriptor_memory_s1            (cpu_instruction_master_granted_descriptor_memory_s1),
      .cpu_instruction_master_granted_ext_flash_s1                    (cpu_instruction_master_granted_ext_flash_s1),
      .cpu_instruction_master_granted_onchip_memory_s1                (cpu_instruction_master_granted_onchip_memory_s1),
      .cpu_instruction_master_latency_counter                         (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_qualified_request_descriptor_memory_s1  (cpu_instruction_master_qualified_request_descriptor_memory_s1),
      .cpu_instruction_master_qualified_request_ext_flash_s1          (cpu_instruction_master_qualified_request_ext_flash_s1),
      .cpu_instruction_master_qualified_request_onchip_memory_s1      (cpu_instruction_master_qualified_request_onchip_memory_s1),
      .cpu_instruction_master_read                                    (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module   (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_descriptor_memory_s1    (cpu_instruction_master_read_data_valid_descriptor_memory_s1),
      .cpu_instruction_master_read_data_valid_ext_flash_s1            (cpu_instruction_master_read_data_valid_ext_flash_s1),
      .cpu_instruction_master_read_data_valid_onchip_memory_s1        (cpu_instruction_master_read_data_valid_onchip_memory_s1),
      .cpu_instruction_master_readdata                                (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                           (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_cpu_jtag_debug_module          (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_instruction_master_requests_descriptor_memory_s1           (cpu_instruction_master_requests_descriptor_memory_s1),
      .cpu_instruction_master_requests_ext_flash_s1                   (cpu_instruction_master_requests_ext_flash_s1),
      .cpu_instruction_master_requests_onchip_memory_s1               (cpu_instruction_master_requests_onchip_memory_s1),
      .cpu_instruction_master_waitrequest                             (cpu_instruction_master_waitrequest),
      .cpu_jtag_debug_module_readdata_from_sa                         (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                              (d1_cpu_jtag_debug_module_end_xfer),
      .d1_descriptor_memory_s1_end_xfer                               (d1_descriptor_memory_s1_end_xfer),
      .d1_flash_tristate_bridge_avalon_slave_end_xfer                 (d1_flash_tristate_bridge_avalon_slave_end_xfer),
      .d1_onchip_memory_s1_end_xfer                                   (d1_onchip_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                          (descriptor_memory_s1_readdata_from_sa),
      .ext_flash_s1_wait_counter_eq_0                                 (ext_flash_s1_wait_counter_eq_0),
      .incoming_flash_tristate_bridge_data                            (incoming_flash_tristate_bridge_data),
      .onchip_memory_s1_readdata_from_sa                              (onchip_memory_s1_readdata_from_sa),
      .reset_n                                                        (pll_sys_clk_reset_n)
    );

  cpu the_cpu
    (
      .clk                                   (pll_sys_clk),
      .d_address                             (cpu_data_master_address),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  ddr2_s1_arbitrator the_ddr2_s1
    (
      .SS_OCT_SOPC_burst_0_downstream_address_to_slave                       (SS_OCT_SOPC_burst_0_downstream_address_to_slave),
      .SS_OCT_SOPC_burst_0_downstream_arbitrationshare                       (SS_OCT_SOPC_burst_0_downstream_arbitrationshare),
      .SS_OCT_SOPC_burst_0_downstream_burstcount                             (SS_OCT_SOPC_burst_0_downstream_burstcount),
      .SS_OCT_SOPC_burst_0_downstream_byteenable                             (SS_OCT_SOPC_burst_0_downstream_byteenable),
      .SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1                        (SS_OCT_SOPC_burst_0_downstream_granted_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_latency_counter                        (SS_OCT_SOPC_burst_0_downstream_latency_counter),
      .SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1              (SS_OCT_SOPC_burst_0_downstream_qualified_request_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_read                                   (SS_OCT_SOPC_burst_0_downstream_read),
      .SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1                (SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register (SS_OCT_SOPC_burst_0_downstream_read_data_valid_ddr2_s1_shift_register),
      .SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1                       (SS_OCT_SOPC_burst_0_downstream_requests_ddr2_s1),
      .SS_OCT_SOPC_burst_0_downstream_write                                  (SS_OCT_SOPC_burst_0_downstream_write),
      .SS_OCT_SOPC_burst_0_downstream_writedata                              (SS_OCT_SOPC_burst_0_downstream_writedata),
      .clk                                                                   (ddr2_phy_clk_out),
      .d1_ddr2_s1_end_xfer                                                   (d1_ddr2_s1_end_xfer),
      .ddr2_s1_address                                                       (ddr2_s1_address),
      .ddr2_s1_beginbursttransfer                                            (ddr2_s1_beginbursttransfer),
      .ddr2_s1_burstcount                                                    (ddr2_s1_burstcount),
      .ddr2_s1_byteenable                                                    (ddr2_s1_byteenable),
      .ddr2_s1_read                                                          (ddr2_s1_read),
      .ddr2_s1_readdata                                                      (ddr2_s1_readdata),
      .ddr2_s1_readdata_from_sa                                              (ddr2_s1_readdata_from_sa),
      .ddr2_s1_readdatavalid                                                 (ddr2_s1_readdatavalid),
      .ddr2_s1_resetrequest_n                                                (ddr2_s1_resetrequest_n),
      .ddr2_s1_resetrequest_n_from_sa                                        (ddr2_s1_resetrequest_n_from_sa),
      .ddr2_s1_waitrequest_n                                                 (ddr2_s1_waitrequest_n),
      .ddr2_s1_waitrequest_n_from_sa                                         (ddr2_s1_waitrequest_n_from_sa),
      .ddr2_s1_write                                                         (ddr2_s1_write),
      .ddr2_s1_writedata                                                     (ddr2_s1_writedata),
      .pipeline_bridge_ddr2_m1_address_to_slave                              (pipeline_bridge_ddr2_m1_address_to_slave),
      .pipeline_bridge_ddr2_m1_burstcount                                    (pipeline_bridge_ddr2_m1_burstcount),
      .pipeline_bridge_ddr2_m1_byteenable                                    (pipeline_bridge_ddr2_m1_byteenable),
      .pipeline_bridge_ddr2_m1_chipselect                                    (pipeline_bridge_ddr2_m1_chipselect),
      .pipeline_bridge_ddr2_m1_granted_ddr2_s1                               (pipeline_bridge_ddr2_m1_granted_ddr2_s1),
      .pipeline_bridge_ddr2_m1_latency_counter                               (pipeline_bridge_ddr2_m1_latency_counter),
      .pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1                     (pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1),
      .pipeline_bridge_ddr2_m1_read                                          (pipeline_bridge_ddr2_m1_read),
      .pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1                       (pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1),
      .pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register        (pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register),
      .pipeline_bridge_ddr2_m1_requests_ddr2_s1                              (pipeline_bridge_ddr2_m1_requests_ddr2_s1),
      .pipeline_bridge_ddr2_m1_write                                         (pipeline_bridge_ddr2_m1_write),
      .pipeline_bridge_ddr2_m1_writedata                                     (pipeline_bridge_ddr2_m1_writedata),
      .reset_n                                                               (ddr2_phy_clk_out_reset_n)
    );

  //ddr2_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr2_aux_full_rate_clk_out = out_clk_ddr2_aux_full_rate_clk;

  //ddr2_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr2_aux_half_rate_clk_out = out_clk_ddr2_aux_half_rate_clk;

  //ddr2_phy_clk_out out_clk assignment, which is an e_assign
  assign ddr2_phy_clk_out = out_clk_ddr2_phy_clk;

  //reset is asserted asynchronously and deasserted synchronously
  SS_OCT_SOPC_reset_clk_50_domain_synch_module SS_OCT_SOPC_reset_clk_50_domain_synch
    (
      .clk      (clk_50),
      .data_in  (1'b1),
      .data_out (clk_50_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa |
    ~ddr2_s1_resetrequest_n_from_sa |
    ~ddr2_s1_resetrequest_n_from_sa |
    pll_s1_resetrequest_from_sa |
    pll_s1_resetrequest_from_sa);

  ddr2 the_ddr2
    (
      .aux_full_rate_clk     (out_clk_ddr2_aux_full_rate_clk),
      .aux_half_rate_clk     (out_clk_ddr2_aux_half_rate_clk),
      .aux_scan_clk          (aux_scan_clk_from_the_ddr2),
      .aux_scan_clk_reset_n  (aux_scan_clk_reset_n_from_the_ddr2),
      .dll_reference_clk     (dll_reference_clk_from_the_ddr2),
      .dqs_delay_ctrl_export (dqs_delay_ctrl_export_from_the_ddr2),
      .global_reset_n        (global_reset_n_to_the_ddr2),
      .local_address         (ddr2_s1_address),
      .local_be              (ddr2_s1_byteenable),
      .local_burstbegin      (ddr2_s1_beginbursttransfer),
      .local_init_done       (local_init_done_from_the_ddr2),
      .local_rdata           (ddr2_s1_readdata),
      .local_rdata_valid     (ddr2_s1_readdatavalid),
      .local_read_req        (ddr2_s1_read),
      .local_ready           (ddr2_s1_waitrequest_n),
      .local_refresh_ack     (local_refresh_ack_from_the_ddr2),
      .local_size            (ddr2_s1_burstcount),
      .local_wdata           (ddr2_s1_writedata),
      .local_wdata_req       (local_wdata_req_from_the_ddr2),
      .local_write_req       (ddr2_s1_write),
      .mem_addr              (mem_addr_from_the_ddr2),
      .mem_ba                (mem_ba_from_the_ddr2),
      .mem_cas_n             (mem_cas_n_from_the_ddr2),
      .mem_cke               (mem_cke_from_the_ddr2),
      .mem_clk               (mem_clk_to_and_from_the_ddr2),
      .mem_clk_n             (mem_clk_n_to_and_from_the_ddr2),
      .mem_cs_n              (mem_cs_n_from_the_ddr2),
      .mem_dm                (mem_dm_from_the_ddr2),
      .mem_dq                (mem_dq_to_and_from_the_ddr2),
      .mem_dqs               (mem_dqs_to_and_from_the_ddr2),
      .mem_dqsn              (mem_dqsn_to_and_from_the_ddr2),
      .mem_odt               (mem_odt_from_the_ddr2),
      .mem_ras_n             (mem_ras_n_from_the_ddr2),
      .mem_we_n              (mem_we_n_from_the_ddr2),
      .oct_ctl_rs_value      (oct_ctl_rs_value_to_the_ddr2),
      .oct_ctl_rt_value      (oct_ctl_rt_value_to_the_ddr2),
      .phy_clk               (out_clk_ddr2_phy_clk),
      .pll_ref_clk           (clk_50),
      .reset_phy_clk_n       (reset_phy_clk_n_from_the_ddr2),
      .reset_request_n       (ddr2_s1_resetrequest_n),
      .soft_reset_n          (clk_50_reset_n)
    );

  descriptor_memory_s1_arbitrator the_descriptor_memory_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_granted_descriptor_memory_s1                              (cpu_data_master_granted_descriptor_memory_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_descriptor_memory_s1                    (cpu_data_master_qualified_request_descriptor_memory_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_descriptor_memory_s1                      (cpu_data_master_read_data_valid_descriptor_memory_s1),
      .cpu_data_master_requests_descriptor_memory_s1                             (cpu_data_master_requests_descriptor_memory_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                   (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_descriptor_memory_s1                       (cpu_instruction_master_granted_descriptor_memory_s1),
      .cpu_instruction_master_latency_counter                                    (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_descriptor_memory_s1             (cpu_instruction_master_qualified_request_descriptor_memory_s1),
      .cpu_instruction_master_read                                               (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_descriptor_memory_s1               (cpu_instruction_master_read_data_valid_descriptor_memory_s1),
      .cpu_instruction_master_requests_descriptor_memory_s1                      (cpu_instruction_master_requests_descriptor_memory_s1),
      .d1_descriptor_memory_s1_end_xfer                                          (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_address                                              (descriptor_memory_s1_address),
      .descriptor_memory_s1_byteenable                                           (descriptor_memory_s1_byteenable),
      .descriptor_memory_s1_chipselect                                           (descriptor_memory_s1_chipselect),
      .descriptor_memory_s1_clken                                                (descriptor_memory_s1_clken),
      .descriptor_memory_s1_readdata                                             (descriptor_memory_s1_readdata),
      .descriptor_memory_s1_readdata_from_sa                                     (descriptor_memory_s1_readdata_from_sa),
      .descriptor_memory_s1_write                                                (descriptor_memory_s1_write),
      .descriptor_memory_s1_writedata                                            (descriptor_memory_s1_writedata),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sgdma_rx_descriptor_read_address_to_slave                                 (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_descriptor_memory_s1                     (sgdma_rx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                                  (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1           (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                             (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1             (sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_requests_descriptor_memory_s1                    (sgdma_rx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_address_to_slave                                (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_descriptor_memory_s1                    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1          (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_descriptor_memory_s1                   (sgdma_rx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_write                                           (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                                       (sgdma_rx_descriptor_write_writedata),
      .sgdma_tx_descriptor_read_address_to_slave                                 (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_descriptor_memory_s1                     (sgdma_tx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                                  (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1           (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                             (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1             (sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_requests_descriptor_memory_s1                    (sgdma_tx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_address_to_slave                                (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_descriptor_memory_s1                    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1          (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_descriptor_memory_s1                   (sgdma_tx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_write                                           (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                                       (sgdma_tx_descriptor_write_writedata)
    );

  descriptor_memory the_descriptor_memory
    (
      .address    (descriptor_memory_s1_address),
      .byteenable (descriptor_memory_s1_byteenable),
      .chipselect (descriptor_memory_s1_chipselect),
      .clk        (pll_sys_clk),
      .clken      (descriptor_memory_s1_clken),
      .readdata   (descriptor_memory_s1_readdata),
      .write      (descriptor_memory_s1_write),
      .writedata  (descriptor_memory_s1_writedata)
    );

  flash_tristate_bridge_avalon_slave_arbitrator the_flash_tristate_bridge_avalon_slave
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_byteenable_ext_flash_s1                                   (cpu_data_master_byteenable_ext_flash_s1),
      .cpu_data_master_dbs_address                                               (cpu_data_master_dbs_address),
      .cpu_data_master_dbs_write_16                                              (cpu_data_master_dbs_write_16),
      .cpu_data_master_granted_ext_flash_s1                                      (cpu_data_master_granted_ext_flash_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_ext_flash_s1                            (cpu_data_master_qualified_request_ext_flash_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_ext_flash_s1                              (cpu_data_master_read_data_valid_ext_flash_s1),
      .cpu_data_master_requests_ext_flash_s1                                     (cpu_data_master_requests_ext_flash_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_instruction_master_address_to_slave                                   (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_dbs_address                                        (cpu_instruction_master_dbs_address),
      .cpu_instruction_master_granted_ext_flash_s1                               (cpu_instruction_master_granted_ext_flash_s1),
      .cpu_instruction_master_latency_counter                                    (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_ext_flash_s1                     (cpu_instruction_master_qualified_request_ext_flash_s1),
      .cpu_instruction_master_read                                               (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_ext_flash_s1                       (cpu_instruction_master_read_data_valid_ext_flash_s1),
      .cpu_instruction_master_requests_ext_flash_s1                              (cpu_instruction_master_requests_ext_flash_s1),
      .d1_flash_tristate_bridge_avalon_slave_end_xfer                            (d1_flash_tristate_bridge_avalon_slave_end_xfer),
      .ext_flash_s1_wait_counter_eq_0                                            (ext_flash_s1_wait_counter_eq_0),
      .flash_tristate_bridge_address                                             (flash_tristate_bridge_address),
      .flash_tristate_bridge_data                                                (flash_tristate_bridge_data),
      .flash_tristate_bridge_readn                                               (flash_tristate_bridge_readn),
      .flash_tristate_bridge_writen                                              (flash_tristate_bridge_writen),
      .incoming_flash_tristate_bridge_data                                       (incoming_flash_tristate_bridge_data),
      .incoming_flash_tristate_bridge_data_with_Xs_converted_to_0                (incoming_flash_tristate_bridge_data_with_Xs_converted_to_0),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .select_n_to_the_ext_flash                                                 (select_n_to_the_ext_flash)
    );

  high_res_timer_s1_arbitrator the_high_res_timer_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_high_res_timer_s1                                 (cpu_data_master_granted_high_res_timer_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_high_res_timer_s1                       (cpu_data_master_qualified_request_high_res_timer_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_high_res_timer_s1                         (cpu_data_master_read_data_valid_high_res_timer_s1),
      .cpu_data_master_requests_high_res_timer_s1                                (cpu_data_master_requests_high_res_timer_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_high_res_timer_s1_end_xfer                                             (d1_high_res_timer_s1_end_xfer),
      .high_res_timer_s1_address                                                 (high_res_timer_s1_address),
      .high_res_timer_s1_chipselect                                              (high_res_timer_s1_chipselect),
      .high_res_timer_s1_irq                                                     (high_res_timer_s1_irq),
      .high_res_timer_s1_irq_from_sa                                             (high_res_timer_s1_irq_from_sa),
      .high_res_timer_s1_readdata                                                (high_res_timer_s1_readdata),
      .high_res_timer_s1_readdata_from_sa                                        (high_res_timer_s1_readdata_from_sa),
      .high_res_timer_s1_reset_n                                                 (high_res_timer_s1_reset_n),
      .high_res_timer_s1_write_n                                                 (high_res_timer_s1_write_n),
      .high_res_timer_s1_writedata                                               (high_res_timer_s1_writedata),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  high_res_timer the_high_res_timer
    (
      .address    (high_res_timer_s1_address),
      .chipselect (high_res_timer_s1_chipselect),
      .clk        (pll_sys_clk),
      .irq        (high_res_timer_s1_irq),
      .readdata   (high_res_timer_s1_readdata),
      .reset_n    (high_res_timer_s1_reset_n),
      .write_n    (high_res_timer_s1_write_n),
      .writedata  (high_res_timer_s1_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_jtag_uart_avalon_jtag_slave                       (cpu_data_master_granted_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave             (cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave               (cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_requests_jtag_uart_avalon_jtag_slave                      (cpu_data_master_requests_jtag_uart_avalon_jtag_slave),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                   (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                                       (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                                    (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                                 (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa                         (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                                           (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                   (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                                        (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                                      (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                              (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                                  (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa                          (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                                       (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                                   (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                           (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                                       (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                                     (jtag_uart_avalon_jtag_slave_writedata),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (pll_sys_clk),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  master_read_avalon_master_arbitrator the_master_read_avalon_master
    (
      .clk                                                                      (clk_50),
      .clock_crossing_master_ddr2_s1_readdata_from_sa                           (clock_crossing_master_ddr2_s1_readdata_from_sa),
      .clock_crossing_master_ddr2_s1_waitrequest_from_sa                        (clock_crossing_master_ddr2_s1_waitrequest_from_sa),
      .d1_clock_crossing_master_ddr2_s1_end_xfer                                (d1_clock_crossing_master_ddr2_s1_end_xfer),
      .master_read_avalon_master_address                                        (master_read_avalon_master_address),
      .master_read_avalon_master_address_to_slave                               (master_read_avalon_master_address_to_slave),
      .master_read_avalon_master_burstcount                                     (master_read_avalon_master_burstcount),
      .master_read_avalon_master_byteenable                                     (master_read_avalon_master_byteenable),
      .master_read_avalon_master_read                                           (master_read_avalon_master_read),
      .master_read_avalon_master_readdata                                       (master_read_avalon_master_readdata),
      .master_read_avalon_master_readdatavalid                                  (master_read_avalon_master_readdatavalid),
      .master_read_avalon_master_reset                                          (master_read_avalon_master_reset),
      .master_read_avalon_master_waitrequest                                    (master_read_avalon_master_waitrequest),
      .master_read_granted_clock_crossing_master_ddr2_s1                        (master_read_granted_clock_crossing_master_ddr2_s1),
      .master_read_latency_counter                                              (master_read_latency_counter),
      .master_read_qualified_request_clock_crossing_master_ddr2_s1              (master_read_qualified_request_clock_crossing_master_ddr2_s1),
      .master_read_read_data_valid_clock_crossing_master_ddr2_s1                (master_read_read_data_valid_clock_crossing_master_ddr2_s1),
      .master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register (master_read_read_data_valid_clock_crossing_master_ddr2_s1_shift_register),
      .master_read_requests_clock_crossing_master_ddr2_s1                       (master_read_requests_clock_crossing_master_ddr2_s1),
      .reset_n                                                                  (clk_50_reset_n)
    );

  master_read the_master_read
    (
      .clk                     (clk_50),
      .control_done            (control_done_from_the_master_read),
      .control_early_done      (control_early_done_from_the_master_read),
      .control_fixed_location  (control_fixed_location_to_the_master_read),
      .control_go              (control_go_to_the_master_read),
      .control_read_base       (control_read_base_to_the_master_read),
      .control_read_length     (control_read_length_to_the_master_read),
      .master_address          (master_read_avalon_master_address),
      .master_burstcount       (master_read_avalon_master_burstcount),
      .master_byteenable       (master_read_avalon_master_byteenable),
      .master_read             (master_read_avalon_master_read),
      .master_readdata         (master_read_avalon_master_readdata),
      .master_readdatavalid    (master_read_avalon_master_readdatavalid),
      .master_waitrequest      (master_read_avalon_master_waitrequest),
      .reset                   (master_read_avalon_master_reset),
      .user_buffer_output_data (user_buffer_output_data_from_the_master_read),
      .user_data_available     (user_data_available_from_the_master_read),
      .user_read_buffer        (user_read_buffer_to_the_master_read)
    );

  master_write_avalon_master_arbitrator the_master_write_avalon_master
    (
      .clk                                                          (clk_50),
      .clock_crossing_master_ddr2_s1_waitrequest_from_sa            (clock_crossing_master_ddr2_s1_waitrequest_from_sa),
      .d1_clock_crossing_master_ddr2_s1_end_xfer                    (d1_clock_crossing_master_ddr2_s1_end_xfer),
      .master_write_avalon_master_address                           (master_write_avalon_master_address),
      .master_write_avalon_master_address_to_slave                  (master_write_avalon_master_address_to_slave),
      .master_write_avalon_master_burstcount                        (master_write_avalon_master_burstcount),
      .master_write_avalon_master_byteenable                        (master_write_avalon_master_byteenable),
      .master_write_avalon_master_reset                             (master_write_avalon_master_reset),
      .master_write_avalon_master_waitrequest                       (master_write_avalon_master_waitrequest),
      .master_write_avalon_master_write                             (master_write_avalon_master_write),
      .master_write_avalon_master_writedata                         (master_write_avalon_master_writedata),
      .master_write_granted_clock_crossing_master_ddr2_s1           (master_write_granted_clock_crossing_master_ddr2_s1),
      .master_write_qualified_request_clock_crossing_master_ddr2_s1 (master_write_qualified_request_clock_crossing_master_ddr2_s1),
      .master_write_requests_clock_crossing_master_ddr2_s1          (master_write_requests_clock_crossing_master_ddr2_s1),
      .reset_n                                                      (clk_50_reset_n)
    );

  master_write the_master_write
    (
      .clk                    (clk_50),
      .control_done           (control_done_from_the_master_write),
      .control_fixed_location (control_fixed_location_to_the_master_write),
      .control_go             (control_go_to_the_master_write),
      .control_write_base     (control_write_base_to_the_master_write),
      .control_write_length   (control_write_length_to_the_master_write),
      .master_address         (master_write_avalon_master_address),
      .master_burstcount      (master_write_avalon_master_burstcount),
      .master_byteenable      (master_write_avalon_master_byteenable),
      .master_waitrequest     (master_write_avalon_master_waitrequest),
      .master_write           (master_write_avalon_master_write),
      .master_writedata       (master_write_avalon_master_writedata),
      .reset                  (master_write_avalon_master_reset),
      .user_buffer_full       (user_buffer_full_from_the_master_write),
      .user_buffer_input_data (user_buffer_input_data_to_the_master_write),
      .user_write_buffer      (user_write_buffer_to_the_master_write)
    );

  onchip_memory_s1_arbitrator the_onchip_memory_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_granted_onchip_memory_s1                                  (cpu_data_master_granted_onchip_memory_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_onchip_memory_s1                        (cpu_data_master_qualified_request_onchip_memory_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_onchip_memory_s1                          (cpu_data_master_read_data_valid_onchip_memory_s1),
      .cpu_data_master_requests_onchip_memory_s1                                 (cpu_data_master_requests_onchip_memory_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                   (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_onchip_memory_s1                           (cpu_instruction_master_granted_onchip_memory_s1),
      .cpu_instruction_master_latency_counter                                    (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_onchip_memory_s1                 (cpu_instruction_master_qualified_request_onchip_memory_s1),
      .cpu_instruction_master_read                                               (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_onchip_memory_s1                   (cpu_instruction_master_read_data_valid_onchip_memory_s1),
      .cpu_instruction_master_requests_onchip_memory_s1                          (cpu_instruction_master_requests_onchip_memory_s1),
      .d1_onchip_memory_s1_end_xfer                                              (d1_onchip_memory_s1_end_xfer),
      .onchip_memory_s1_address                                                  (onchip_memory_s1_address),
      .onchip_memory_s1_byteenable                                               (onchip_memory_s1_byteenable),
      .onchip_memory_s1_chipselect                                               (onchip_memory_s1_chipselect),
      .onchip_memory_s1_clken                                                    (onchip_memory_s1_clken),
      .onchip_memory_s1_readdata                                                 (onchip_memory_s1_readdata),
      .onchip_memory_s1_readdata_from_sa                                         (onchip_memory_s1_readdata_from_sa),
      .onchip_memory_s1_write                                                    (onchip_memory_s1_write),
      .onchip_memory_s1_writedata                                                (onchip_memory_s1_writedata),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sgdma_rx_m_write_address_to_slave                                         (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                                               (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_onchip_memory_s1                                 (sgdma_rx_m_write_granted_onchip_memory_s1),
      .sgdma_rx_m_write_qualified_request_onchip_memory_s1                       (sgdma_rx_m_write_qualified_request_onchip_memory_s1),
      .sgdma_rx_m_write_requests_onchip_memory_s1                                (sgdma_rx_m_write_requests_onchip_memory_s1),
      .sgdma_rx_m_write_write                                                    (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                                                (sgdma_rx_m_write_writedata),
      .sgdma_tx_m_read_address_to_slave                                          (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_onchip_memory_s1                                  (sgdma_tx_m_read_granted_onchip_memory_s1),
      .sgdma_tx_m_read_latency_counter                                           (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_onchip_memory_s1                        (sgdma_tx_m_read_qualified_request_onchip_memory_s1),
      .sgdma_tx_m_read_read                                                      (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_onchip_memory_s1                          (sgdma_tx_m_read_read_data_valid_onchip_memory_s1),
      .sgdma_tx_m_read_requests_onchip_memory_s1                                 (sgdma_tx_m_read_requests_onchip_memory_s1)
    );

  onchip_memory the_onchip_memory
    (
      .address    (onchip_memory_s1_address),
      .byteenable (onchip_memory_s1_byteenable),
      .chipselect (onchip_memory_s1_chipselect),
      .clk        (pll_sys_clk),
      .clken      (onchip_memory_s1_clken),
      .readdata   (onchip_memory_s1_readdata),
      .write      (onchip_memory_s1_write),
      .writedata  (onchip_memory_s1_writedata)
    );

  packet_memory_s1_arbitrator the_packet_memory_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                (cpu_data_master_byteenable),
      .cpu_data_master_granted_packet_memory_s1                                  (cpu_data_master_granted_packet_memory_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_packet_memory_s1                        (cpu_data_master_qualified_request_packet_memory_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_packet_memory_s1                          (cpu_data_master_read_data_valid_packet_memory_s1),
      .cpu_data_master_requests_packet_memory_s1                                 (cpu_data_master_requests_packet_memory_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_packet_memory_s1_end_xfer                                              (d1_packet_memory_s1_end_xfer),
      .packet_memory_s1_address                                                  (packet_memory_s1_address),
      .packet_memory_s1_byteenable                                               (packet_memory_s1_byteenable),
      .packet_memory_s1_chipselect                                               (packet_memory_s1_chipselect),
      .packet_memory_s1_clken                                                    (packet_memory_s1_clken),
      .packet_memory_s1_readdata                                                 (packet_memory_s1_readdata),
      .packet_memory_s1_readdata_from_sa                                         (packet_memory_s1_readdata_from_sa),
      .packet_memory_s1_write                                                    (packet_memory_s1_write),
      .packet_memory_s1_writedata                                                (packet_memory_s1_writedata),
      .reset_n                                                                   (pll_sys_clk_reset_n)
    );

  packet_memory_s2_arbitrator the_packet_memory_s2
    (
      .clk                                                 (pll_sys_clk),
      .d1_packet_memory_s2_end_xfer                        (d1_packet_memory_s2_end_xfer),
      .packet_memory_s2_address                            (packet_memory_s2_address),
      .packet_memory_s2_byteenable                         (packet_memory_s2_byteenable),
      .packet_memory_s2_chipselect                         (packet_memory_s2_chipselect),
      .packet_memory_s2_clken                              (packet_memory_s2_clken),
      .packet_memory_s2_readdata                           (packet_memory_s2_readdata),
      .packet_memory_s2_readdata_from_sa                   (packet_memory_s2_readdata_from_sa),
      .packet_memory_s2_write                              (packet_memory_s2_write),
      .packet_memory_s2_writedata                          (packet_memory_s2_writedata),
      .reset_n                                             (pll_sys_clk_reset_n),
      .sgdma_rx_m_write_address_to_slave                   (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                         (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_packet_memory_s2           (sgdma_rx_m_write_granted_packet_memory_s2),
      .sgdma_rx_m_write_qualified_request_packet_memory_s2 (sgdma_rx_m_write_qualified_request_packet_memory_s2),
      .sgdma_rx_m_write_requests_packet_memory_s2          (sgdma_rx_m_write_requests_packet_memory_s2),
      .sgdma_rx_m_write_write                              (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                          (sgdma_rx_m_write_writedata),
      .sgdma_tx_m_read_address_to_slave                    (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_packet_memory_s2            (sgdma_tx_m_read_granted_packet_memory_s2),
      .sgdma_tx_m_read_latency_counter                     (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_packet_memory_s2  (sgdma_tx_m_read_qualified_request_packet_memory_s2),
      .sgdma_tx_m_read_read                                (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_packet_memory_s2    (sgdma_tx_m_read_read_data_valid_packet_memory_s2),
      .sgdma_tx_m_read_requests_packet_memory_s2           (sgdma_tx_m_read_requests_packet_memory_s2)
    );

  packet_memory the_packet_memory
    (
      .address     (packet_memory_s1_address),
      .address2    (packet_memory_s2_address),
      .byteenable  (packet_memory_s1_byteenable),
      .byteenable2 (packet_memory_s2_byteenable),
      .chipselect  (packet_memory_s1_chipselect),
      .chipselect2 (packet_memory_s2_chipselect),
      .clk         (pll_sys_clk),
      .clk2        (pll_sys_clk),
      .clken       (packet_memory_s1_clken),
      .clken2      (packet_memory_s2_clken),
      .readdata    (packet_memory_s1_readdata),
      .readdata2   (packet_memory_s2_readdata),
      .write       (packet_memory_s1_write),
      .write2      (packet_memory_s2_write),
      .writedata   (packet_memory_s1_writedata),
      .writedata2  (packet_memory_s2_writedata)
    );

  pipeline_bridge_ddr2_s1_arbitrator the_pipeline_bridge_ddr2_s1
    (
      .clk                                                                               (ddr2_phy_clk_out),
      .clock_crossing_ddr2_cpu_m1_address_to_slave                                       (clock_crossing_ddr2_cpu_m1_address_to_slave),
      .clock_crossing_ddr2_cpu_m1_byteenable                                             (clock_crossing_ddr2_cpu_m1_byteenable),
      .clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1                        (clock_crossing_ddr2_cpu_m1_granted_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_latency_counter                                        (clock_crossing_ddr2_cpu_m1_latency_counter),
      .clock_crossing_ddr2_cpu_m1_nativeaddress                                          (clock_crossing_ddr2_cpu_m1_nativeaddress),
      .clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1              (clock_crossing_ddr2_cpu_m1_qualified_request_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_read                                                   (clock_crossing_ddr2_cpu_m1_read),
      .clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1                (clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register (clock_crossing_ddr2_cpu_m1_read_data_valid_pipeline_bridge_ddr2_s1_shift_register),
      .clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1                       (clock_crossing_ddr2_cpu_m1_requests_pipeline_bridge_ddr2_s1),
      .clock_crossing_ddr2_cpu_m1_write                                                  (clock_crossing_ddr2_cpu_m1_write),
      .clock_crossing_ddr2_cpu_m1_writedata                                              (clock_crossing_ddr2_cpu_m1_writedata),
      .d1_pipeline_bridge_ddr2_s1_end_xfer                                               (d1_pipeline_bridge_ddr2_s1_end_xfer),
      .pipeline_bridge_ddr2_s1_address                                                   (pipeline_bridge_ddr2_s1_address),
      .pipeline_bridge_ddr2_s1_arbiterlock                                               (pipeline_bridge_ddr2_s1_arbiterlock),
      .pipeline_bridge_ddr2_s1_arbiterlock2                                              (pipeline_bridge_ddr2_s1_arbiterlock2),
      .pipeline_bridge_ddr2_s1_burstcount                                                (pipeline_bridge_ddr2_s1_burstcount),
      .pipeline_bridge_ddr2_s1_byteenable                                                (pipeline_bridge_ddr2_s1_byteenable),
      .pipeline_bridge_ddr2_s1_chipselect                                                (pipeline_bridge_ddr2_s1_chipselect),
      .pipeline_bridge_ddr2_s1_debugaccess                                               (pipeline_bridge_ddr2_s1_debugaccess),
      .pipeline_bridge_ddr2_s1_endofpacket                                               (pipeline_bridge_ddr2_s1_endofpacket),
      .pipeline_bridge_ddr2_s1_endofpacket_from_sa                                       (pipeline_bridge_ddr2_s1_endofpacket_from_sa),
      .pipeline_bridge_ddr2_s1_nativeaddress                                             (pipeline_bridge_ddr2_s1_nativeaddress),
      .pipeline_bridge_ddr2_s1_read                                                      (pipeline_bridge_ddr2_s1_read),
      .pipeline_bridge_ddr2_s1_readdata                                                  (pipeline_bridge_ddr2_s1_readdata),
      .pipeline_bridge_ddr2_s1_readdata_from_sa                                          (pipeline_bridge_ddr2_s1_readdata_from_sa),
      .pipeline_bridge_ddr2_s1_readdatavalid                                             (pipeline_bridge_ddr2_s1_readdatavalid),
      .pipeline_bridge_ddr2_s1_reset_n                                                   (pipeline_bridge_ddr2_s1_reset_n),
      .pipeline_bridge_ddr2_s1_waitrequest                                               (pipeline_bridge_ddr2_s1_waitrequest),
      .pipeline_bridge_ddr2_s1_waitrequest_from_sa                                       (pipeline_bridge_ddr2_s1_waitrequest_from_sa),
      .pipeline_bridge_ddr2_s1_write                                                     (pipeline_bridge_ddr2_s1_write),
      .pipeline_bridge_ddr2_s1_writedata                                                 (pipeline_bridge_ddr2_s1_writedata),
      .reset_n                                                                           (ddr2_phy_clk_out_reset_n)
    );

  pipeline_bridge_ddr2_m1_arbitrator the_pipeline_bridge_ddr2_m1
    (
      .clk                                                            (ddr2_phy_clk_out),
      .d1_ddr2_s1_end_xfer                                            (d1_ddr2_s1_end_xfer),
      .ddr2_s1_readdata_from_sa                                       (ddr2_s1_readdata_from_sa),
      .ddr2_s1_waitrequest_n_from_sa                                  (ddr2_s1_waitrequest_n_from_sa),
      .pipeline_bridge_ddr2_m1_address                                (pipeline_bridge_ddr2_m1_address),
      .pipeline_bridge_ddr2_m1_address_to_slave                       (pipeline_bridge_ddr2_m1_address_to_slave),
      .pipeline_bridge_ddr2_m1_burstcount                             (pipeline_bridge_ddr2_m1_burstcount),
      .pipeline_bridge_ddr2_m1_byteenable                             (pipeline_bridge_ddr2_m1_byteenable),
      .pipeline_bridge_ddr2_m1_chipselect                             (pipeline_bridge_ddr2_m1_chipselect),
      .pipeline_bridge_ddr2_m1_granted_ddr2_s1                        (pipeline_bridge_ddr2_m1_granted_ddr2_s1),
      .pipeline_bridge_ddr2_m1_latency_counter                        (pipeline_bridge_ddr2_m1_latency_counter),
      .pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1              (pipeline_bridge_ddr2_m1_qualified_request_ddr2_s1),
      .pipeline_bridge_ddr2_m1_read                                   (pipeline_bridge_ddr2_m1_read),
      .pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1                (pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1),
      .pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register (pipeline_bridge_ddr2_m1_read_data_valid_ddr2_s1_shift_register),
      .pipeline_bridge_ddr2_m1_readdata                               (pipeline_bridge_ddr2_m1_readdata),
      .pipeline_bridge_ddr2_m1_readdatavalid                          (pipeline_bridge_ddr2_m1_readdatavalid),
      .pipeline_bridge_ddr2_m1_requests_ddr2_s1                       (pipeline_bridge_ddr2_m1_requests_ddr2_s1),
      .pipeline_bridge_ddr2_m1_waitrequest                            (pipeline_bridge_ddr2_m1_waitrequest),
      .pipeline_bridge_ddr2_m1_write                                  (pipeline_bridge_ddr2_m1_write),
      .pipeline_bridge_ddr2_m1_writedata                              (pipeline_bridge_ddr2_m1_writedata),
      .reset_n                                                        (ddr2_phy_clk_out_reset_n)
    );

  pipeline_bridge_ddr2 the_pipeline_bridge_ddr2
    (
      .clk              (ddr2_phy_clk_out),
      .m1_address       (pipeline_bridge_ddr2_m1_address),
      .m1_burstcount    (pipeline_bridge_ddr2_m1_burstcount),
      .m1_byteenable    (pipeline_bridge_ddr2_m1_byteenable),
      .m1_chipselect    (pipeline_bridge_ddr2_m1_chipselect),
      .m1_debugaccess   (pipeline_bridge_ddr2_m1_debugaccess),
      .m1_endofpacket   (pipeline_bridge_ddr2_m1_endofpacket),
      .m1_read          (pipeline_bridge_ddr2_m1_read),
      .m1_readdata      (pipeline_bridge_ddr2_m1_readdata),
      .m1_readdatavalid (pipeline_bridge_ddr2_m1_readdatavalid),
      .m1_waitrequest   (pipeline_bridge_ddr2_m1_waitrequest),
      .m1_write         (pipeline_bridge_ddr2_m1_write),
      .m1_writedata     (pipeline_bridge_ddr2_m1_writedata),
      .reset_n          (pipeline_bridge_ddr2_s1_reset_n),
      .s1_address       (pipeline_bridge_ddr2_s1_address),
      .s1_arbiterlock   (pipeline_bridge_ddr2_s1_arbiterlock),
      .s1_arbiterlock2  (pipeline_bridge_ddr2_s1_arbiterlock2),
      .s1_burstcount    (pipeline_bridge_ddr2_s1_burstcount),
      .s1_byteenable    (pipeline_bridge_ddr2_s1_byteenable),
      .s1_chipselect    (pipeline_bridge_ddr2_s1_chipselect),
      .s1_debugaccess   (pipeline_bridge_ddr2_s1_debugaccess),
      .s1_endofpacket   (pipeline_bridge_ddr2_s1_endofpacket),
      .s1_nativeaddress (pipeline_bridge_ddr2_s1_nativeaddress),
      .s1_read          (pipeline_bridge_ddr2_s1_read),
      .s1_readdata      (pipeline_bridge_ddr2_s1_readdata),
      .s1_readdatavalid (pipeline_bridge_ddr2_s1_readdatavalid),
      .s1_waitrequest   (pipeline_bridge_ddr2_s1_waitrequest),
      .s1_write         (pipeline_bridge_ddr2_s1_write),
      .s1_writedata     (pipeline_bridge_ddr2_s1_writedata)
    );

  pll_s1_arbitrator the_pll_s1
    (
      .SS_OCT_SOPC_clock_0_out_address_to_slave         (SS_OCT_SOPC_clock_0_out_address_to_slave),
      .SS_OCT_SOPC_clock_0_out_granted_pll_s1           (SS_OCT_SOPC_clock_0_out_granted_pll_s1),
      .SS_OCT_SOPC_clock_0_out_nativeaddress            (SS_OCT_SOPC_clock_0_out_nativeaddress),
      .SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1 (SS_OCT_SOPC_clock_0_out_qualified_request_pll_s1),
      .SS_OCT_SOPC_clock_0_out_read                     (SS_OCT_SOPC_clock_0_out_read),
      .SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1   (SS_OCT_SOPC_clock_0_out_read_data_valid_pll_s1),
      .SS_OCT_SOPC_clock_0_out_requests_pll_s1          (SS_OCT_SOPC_clock_0_out_requests_pll_s1),
      .SS_OCT_SOPC_clock_0_out_write                    (SS_OCT_SOPC_clock_0_out_write),
      .SS_OCT_SOPC_clock_0_out_writedata                (SS_OCT_SOPC_clock_0_out_writedata),
      .clk                                              (clk_50),
      .d1_pll_s1_end_xfer                               (d1_pll_s1_end_xfer),
      .pll_s1_address                                   (pll_s1_address),
      .pll_s1_chipselect                                (pll_s1_chipselect),
      .pll_s1_read                                      (pll_s1_read),
      .pll_s1_readdata                                  (pll_s1_readdata),
      .pll_s1_readdata_from_sa                          (pll_s1_readdata_from_sa),
      .pll_s1_reset_n                                   (pll_s1_reset_n),
      .pll_s1_resetrequest                              (pll_s1_resetrequest),
      .pll_s1_resetrequest_from_sa                      (pll_s1_resetrequest_from_sa),
      .pll_s1_write                                     (pll_s1_write),
      .pll_s1_writedata                                 (pll_s1_writedata),
      .reset_n                                          (clk_50_reset_n)
    );

  //pll_sys_clk out_clk assignment, which is an e_assign
  assign pll_sys_clk = out_clk_pll_c0;

  pll the_pll
    (
      .address      (pll_s1_address),
      .c0           (out_clk_pll_c0),
      .chipselect   (pll_s1_chipselect),
      .clk          (clk_50),
      .read         (pll_s1_read),
      .readdata     (pll_s1_readdata),
      .reset_n      (pll_s1_reset_n),
      .resetrequest (pll_s1_resetrequest),
      .write        (pll_s1_write),
      .writedata    (pll_s1_writedata)
    );

  sgdma_rx_csr_arbitrator the_sgdma_rx_csr
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sgdma_rx_csr                                      (cpu_data_master_granted_sgdma_rx_csr),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sgdma_rx_csr                            (cpu_data_master_qualified_request_sgdma_rx_csr),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_sgdma_rx_csr                              (cpu_data_master_read_data_valid_sgdma_rx_csr),
      .cpu_data_master_requests_sgdma_rx_csr                                     (cpu_data_master_requests_sgdma_rx_csr),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_sgdma_rx_csr_end_xfer                                                  (d1_sgdma_rx_csr_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sgdma_rx_csr_address                                                      (sgdma_rx_csr_address),
      .sgdma_rx_csr_chipselect                                                   (sgdma_rx_csr_chipselect),
      .sgdma_rx_csr_irq                                                          (sgdma_rx_csr_irq),
      .sgdma_rx_csr_irq_from_sa                                                  (sgdma_rx_csr_irq_from_sa),
      .sgdma_rx_csr_read                                                         (sgdma_rx_csr_read),
      .sgdma_rx_csr_readdata                                                     (sgdma_rx_csr_readdata),
      .sgdma_rx_csr_readdata_from_sa                                             (sgdma_rx_csr_readdata_from_sa),
      .sgdma_rx_csr_reset_n                                                      (sgdma_rx_csr_reset_n),
      .sgdma_rx_csr_write                                                        (sgdma_rx_csr_write),
      .sgdma_rx_csr_writedata                                                    (sgdma_rx_csr_writedata)
    );

  sgdma_rx_in_arbitrator the_sgdma_rx_in
    (
      .clk                           (pll_sys_clk),
      .reset_n                       (pll_sys_clk_reset_n),
      .sgdma_rx_in_data              (sgdma_rx_in_data),
      .sgdma_rx_in_empty             (sgdma_rx_in_empty),
      .sgdma_rx_in_endofpacket       (sgdma_rx_in_endofpacket),
      .sgdma_rx_in_error             (sgdma_rx_in_error),
      .sgdma_rx_in_ready             (sgdma_rx_in_ready),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .sgdma_rx_in_startofpacket     (sgdma_rx_in_startofpacket),
      .sgdma_rx_in_valid             (sgdma_rx_in_valid),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  sgdma_rx_descriptor_read_arbitrator the_sgdma_rx_descriptor_read
    (
      .clk                                                             (pll_sys_clk),
      .d1_descriptor_memory_s1_end_xfer                                (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                           (descriptor_memory_s1_readdata_from_sa),
      .reset_n                                                         (pll_sys_clk_reset_n),
      .sgdma_rx_descriptor_read_address                                (sgdma_rx_descriptor_read_address),
      .sgdma_rx_descriptor_read_address_to_slave                       (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_descriptor_memory_s1           (sgdma_rx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                        (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                   (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1   (sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_readdata                               (sgdma_rx_descriptor_read_readdata),
      .sgdma_rx_descriptor_read_readdatavalid                          (sgdma_rx_descriptor_read_readdatavalid),
      .sgdma_rx_descriptor_read_requests_descriptor_memory_s1          (sgdma_rx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_waitrequest                            (sgdma_rx_descriptor_read_waitrequest)
    );

  sgdma_rx_descriptor_write_arbitrator the_sgdma_rx_descriptor_write
    (
      .clk                                                              (pll_sys_clk),
      .d1_descriptor_memory_s1_end_xfer                                 (d1_descriptor_memory_s1_end_xfer),
      .reset_n                                                          (pll_sys_clk_reset_n),
      .sgdma_rx_descriptor_write_address                                (sgdma_rx_descriptor_write_address),
      .sgdma_rx_descriptor_write_address_to_slave                       (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_descriptor_memory_s1           (sgdma_rx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_descriptor_memory_s1          (sgdma_rx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_waitrequest                            (sgdma_rx_descriptor_write_waitrequest),
      .sgdma_rx_descriptor_write_write                                  (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                              (sgdma_rx_descriptor_write_writedata)
    );

  sgdma_rx_m_write_arbitrator the_sgdma_rx_m_write
    (
      .clk                                                 (pll_sys_clk),
      .d1_onchip_memory_s1_end_xfer                        (d1_onchip_memory_s1_end_xfer),
      .d1_packet_memory_s2_end_xfer                        (d1_packet_memory_s2_end_xfer),
      .reset_n                                             (pll_sys_clk_reset_n),
      .sgdma_rx_m_write_address                            (sgdma_rx_m_write_address),
      .sgdma_rx_m_write_address_to_slave                   (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                         (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_onchip_memory_s1           (sgdma_rx_m_write_granted_onchip_memory_s1),
      .sgdma_rx_m_write_granted_packet_memory_s2           (sgdma_rx_m_write_granted_packet_memory_s2),
      .sgdma_rx_m_write_qualified_request_onchip_memory_s1 (sgdma_rx_m_write_qualified_request_onchip_memory_s1),
      .sgdma_rx_m_write_qualified_request_packet_memory_s2 (sgdma_rx_m_write_qualified_request_packet_memory_s2),
      .sgdma_rx_m_write_requests_onchip_memory_s1          (sgdma_rx_m_write_requests_onchip_memory_s1),
      .sgdma_rx_m_write_requests_packet_memory_s2          (sgdma_rx_m_write_requests_packet_memory_s2),
      .sgdma_rx_m_write_waitrequest                        (sgdma_rx_m_write_waitrequest),
      .sgdma_rx_m_write_write                              (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                          (sgdma_rx_m_write_writedata)
    );

  sgdma_rx the_sgdma_rx
    (
      .clk                           (pll_sys_clk),
      .csr_address                   (sgdma_rx_csr_address),
      .csr_chipselect                (sgdma_rx_csr_chipselect),
      .csr_irq                       (sgdma_rx_csr_irq),
      .csr_read                      (sgdma_rx_csr_read),
      .csr_readdata                  (sgdma_rx_csr_readdata),
      .csr_write                     (sgdma_rx_csr_write),
      .csr_writedata                 (sgdma_rx_csr_writedata),
      .descriptor_read_address       (sgdma_rx_descriptor_read_address),
      .descriptor_read_read          (sgdma_rx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_rx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_rx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),
      .in_data                       (sgdma_rx_in_data),
      .in_empty                      (sgdma_rx_in_empty),
      .in_endofpacket                (sgdma_rx_in_endofpacket),
      .in_error                      (sgdma_rx_in_error),
      .in_ready                      (sgdma_rx_in_ready),
      .in_startofpacket              (sgdma_rx_in_startofpacket),
      .in_valid                      (sgdma_rx_in_valid),
      .m_write_address               (sgdma_rx_m_write_address),
      .m_write_byteenable            (sgdma_rx_m_write_byteenable),
      .m_write_waitrequest           (sgdma_rx_m_write_waitrequest),
      .m_write_write                 (sgdma_rx_m_write_write),
      .m_write_writedata             (sgdma_rx_m_write_writedata),
      .system_reset_n                (sgdma_rx_csr_reset_n)
    );

  sgdma_tx_csr_arbitrator the_sgdma_tx_csr
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sgdma_tx_csr                                      (cpu_data_master_granted_sgdma_tx_csr),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sgdma_tx_csr                            (cpu_data_master_qualified_request_sgdma_tx_csr),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_sgdma_tx_csr                              (cpu_data_master_read_data_valid_sgdma_tx_csr),
      .cpu_data_master_requests_sgdma_tx_csr                                     (cpu_data_master_requests_sgdma_tx_csr),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_sgdma_tx_csr_end_xfer                                                  (d1_sgdma_tx_csr_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sgdma_tx_csr_address                                                      (sgdma_tx_csr_address),
      .sgdma_tx_csr_chipselect                                                   (sgdma_tx_csr_chipselect),
      .sgdma_tx_csr_irq                                                          (sgdma_tx_csr_irq),
      .sgdma_tx_csr_irq_from_sa                                                  (sgdma_tx_csr_irq_from_sa),
      .sgdma_tx_csr_read                                                         (sgdma_tx_csr_read),
      .sgdma_tx_csr_readdata                                                     (sgdma_tx_csr_readdata),
      .sgdma_tx_csr_readdata_from_sa                                             (sgdma_tx_csr_readdata_from_sa),
      .sgdma_tx_csr_reset_n                                                      (sgdma_tx_csr_reset_n),
      .sgdma_tx_csr_write                                                        (sgdma_tx_csr_write),
      .sgdma_tx_csr_writedata                                                    (sgdma_tx_csr_writedata)
    );

  sgdma_tx_descriptor_read_arbitrator the_sgdma_tx_descriptor_read
    (
      .clk                                                             (pll_sys_clk),
      .d1_descriptor_memory_s1_end_xfer                                (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                           (descriptor_memory_s1_readdata_from_sa),
      .reset_n                                                         (pll_sys_clk_reset_n),
      .sgdma_tx_descriptor_read_address                                (sgdma_tx_descriptor_read_address),
      .sgdma_tx_descriptor_read_address_to_slave                       (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_descriptor_memory_s1           (sgdma_tx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                        (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                   (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1   (sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_readdata                               (sgdma_tx_descriptor_read_readdata),
      .sgdma_tx_descriptor_read_readdatavalid                          (sgdma_tx_descriptor_read_readdatavalid),
      .sgdma_tx_descriptor_read_requests_descriptor_memory_s1          (sgdma_tx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_waitrequest                            (sgdma_tx_descriptor_read_waitrequest)
    );

  sgdma_tx_descriptor_write_arbitrator the_sgdma_tx_descriptor_write
    (
      .clk                                                              (pll_sys_clk),
      .d1_descriptor_memory_s1_end_xfer                                 (d1_descriptor_memory_s1_end_xfer),
      .reset_n                                                          (pll_sys_clk_reset_n),
      .sgdma_tx_descriptor_write_address                                (sgdma_tx_descriptor_write_address),
      .sgdma_tx_descriptor_write_address_to_slave                       (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_descriptor_memory_s1           (sgdma_tx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_descriptor_memory_s1          (sgdma_tx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_waitrequest                            (sgdma_tx_descriptor_write_waitrequest),
      .sgdma_tx_descriptor_write_write                                  (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                              (sgdma_tx_descriptor_write_writedata)
    );

  sgdma_tx_m_read_arbitrator the_sgdma_tx_m_read
    (
      .clk                                                (pll_sys_clk),
      .d1_onchip_memory_s1_end_xfer                       (d1_onchip_memory_s1_end_xfer),
      .d1_packet_memory_s2_end_xfer                       (d1_packet_memory_s2_end_xfer),
      .onchip_memory_s1_readdata_from_sa                  (onchip_memory_s1_readdata_from_sa),
      .packet_memory_s2_readdata_from_sa                  (packet_memory_s2_readdata_from_sa),
      .reset_n                                            (pll_sys_clk_reset_n),
      .sgdma_tx_m_read_address                            (sgdma_tx_m_read_address),
      .sgdma_tx_m_read_address_to_slave                   (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_onchip_memory_s1           (sgdma_tx_m_read_granted_onchip_memory_s1),
      .sgdma_tx_m_read_granted_packet_memory_s2           (sgdma_tx_m_read_granted_packet_memory_s2),
      .sgdma_tx_m_read_latency_counter                    (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_onchip_memory_s1 (sgdma_tx_m_read_qualified_request_onchip_memory_s1),
      .sgdma_tx_m_read_qualified_request_packet_memory_s2 (sgdma_tx_m_read_qualified_request_packet_memory_s2),
      .sgdma_tx_m_read_read                               (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_onchip_memory_s1   (sgdma_tx_m_read_read_data_valid_onchip_memory_s1),
      .sgdma_tx_m_read_read_data_valid_packet_memory_s2   (sgdma_tx_m_read_read_data_valid_packet_memory_s2),
      .sgdma_tx_m_read_readdata                           (sgdma_tx_m_read_readdata),
      .sgdma_tx_m_read_readdatavalid                      (sgdma_tx_m_read_readdatavalid),
      .sgdma_tx_m_read_requests_onchip_memory_s1          (sgdma_tx_m_read_requests_onchip_memory_s1),
      .sgdma_tx_m_read_requests_packet_memory_s2          (sgdma_tx_m_read_requests_packet_memory_s2),
      .sgdma_tx_m_read_waitrequest                        (sgdma_tx_m_read_waitrequest)
    );

  sgdma_tx_out_arbitrator the_sgdma_tx_out
    (
      .clk                            (pll_sys_clk),
      .reset_n                        (pll_sys_clk_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_ready             (sgdma_tx_out_ready),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa)
    );

  sgdma_tx the_sgdma_tx
    (
      .clk                           (pll_sys_clk),
      .csr_address                   (sgdma_tx_csr_address),
      .csr_chipselect                (sgdma_tx_csr_chipselect),
      .csr_irq                       (sgdma_tx_csr_irq),
      .csr_read                      (sgdma_tx_csr_read),
      .csr_readdata                  (sgdma_tx_csr_readdata),
      .csr_write                     (sgdma_tx_csr_write),
      .csr_writedata                 (sgdma_tx_csr_writedata),
      .descriptor_read_address       (sgdma_tx_descriptor_read_address),
      .descriptor_read_read          (sgdma_tx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_tx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_tx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),
      .m_read_address                (sgdma_tx_m_read_address),
      .m_read_read                   (sgdma_tx_m_read_read),
      .m_read_readdata               (sgdma_tx_m_read_readdata),
      .m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),
      .m_read_waitrequest            (sgdma_tx_m_read_waitrequest),
      .out_data                      (sgdma_tx_out_data),
      .out_empty                     (sgdma_tx_out_empty),
      .out_endofpacket               (sgdma_tx_out_endofpacket),
      .out_error                     (sgdma_tx_out_error),
      .out_ready                     (sgdma_tx_out_ready),
      .out_startofpacket             (sgdma_tx_out_startofpacket),
      .out_valid                     (sgdma_tx_out_valid),
      .system_reset_n                (sgdma_tx_csr_reset_n)
    );

  sys_timer_s1_arbitrator the_sys_timer_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sys_timer_s1                                      (cpu_data_master_granted_sys_timer_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sys_timer_s1                            (cpu_data_master_qualified_request_sys_timer_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_sys_timer_s1                              (cpu_data_master_read_data_valid_sys_timer_s1),
      .cpu_data_master_requests_sys_timer_s1                                     (cpu_data_master_requests_sys_timer_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_sys_timer_s1_end_xfer                                                  (d1_sys_timer_s1_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sys_timer_s1_address                                                      (sys_timer_s1_address),
      .sys_timer_s1_chipselect                                                   (sys_timer_s1_chipselect),
      .sys_timer_s1_irq                                                          (sys_timer_s1_irq),
      .sys_timer_s1_irq_from_sa                                                  (sys_timer_s1_irq_from_sa),
      .sys_timer_s1_readdata                                                     (sys_timer_s1_readdata),
      .sys_timer_s1_readdata_from_sa                                             (sys_timer_s1_readdata_from_sa),
      .sys_timer_s1_reset_n                                                      (sys_timer_s1_reset_n),
      .sys_timer_s1_write_n                                                      (sys_timer_s1_write_n),
      .sys_timer_s1_writedata                                                    (sys_timer_s1_writedata)
    );

  sys_timer the_sys_timer
    (
      .address    (sys_timer_s1_address),
      .chipselect (sys_timer_s1_chipselect),
      .clk        (pll_sys_clk),
      .irq        (sys_timer_s1_irq),
      .readdata   (sys_timer_s1_readdata),
      .reset_n    (sys_timer_s1_reset_n),
      .write_n    (sys_timer_s1_write_n),
      .writedata  (sys_timer_s1_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sysid_control_slave                               (cpu_data_master_granted_sysid_control_slave),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sysid_control_slave                     (cpu_data_master_qualified_request_sysid_control_slave),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_sysid_control_slave                       (cpu_data_master_read_data_valid_sysid_control_slave),
      .cpu_data_master_requests_sysid_control_slave                              (cpu_data_master_requests_sysid_control_slave),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .d1_sysid_control_slave_end_xfer                                           (d1_sysid_control_slave_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .sysid_control_slave_address                                               (sysid_control_slave_address),
      .sysid_control_slave_readdata                                              (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                                      (sysid_control_slave_readdata_from_sa)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .readdata (sysid_control_slave_readdata)
    );

  tse_mac_control_port_arbitrator the_tse_mac_control_port
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_tse_mac_control_port                              (cpu_data_master_granted_tse_mac_control_port),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_tse_mac_control_port                    (cpu_data_master_qualified_request_tse_mac_control_port),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_tse_mac_control_port                      (cpu_data_master_read_data_valid_tse_mac_control_port),
      .cpu_data_master_requests_tse_mac_control_port                             (cpu_data_master_requests_tse_mac_control_port),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_tse_mac_control_port_end_xfer                                          (d1_tse_mac_control_port_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .tse_mac_control_port_address                                              (tse_mac_control_port_address),
      .tse_mac_control_port_read                                                 (tse_mac_control_port_read),
      .tse_mac_control_port_readdata                                             (tse_mac_control_port_readdata),
      .tse_mac_control_port_readdata_from_sa                                     (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_reset                                                (tse_mac_control_port_reset),
      .tse_mac_control_port_waitrequest                                          (tse_mac_control_port_waitrequest),
      .tse_mac_control_port_waitrequest_from_sa                                  (tse_mac_control_port_waitrequest_from_sa),
      .tse_mac_control_port_write                                                (tse_mac_control_port_write),
      .tse_mac_control_port_writedata                                            (tse_mac_control_port_writedata)
    );

  tse_mac_transmit_arbitrator the_tse_mac_transmit
    (
      .clk                            (pll_sys_clk),
      .reset_n                        (pll_sys_clk_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_data          (tse_mac_transmit_data),
      .tse_mac_transmit_empty         (tse_mac_transmit_empty),
      .tse_mac_transmit_endofpacket   (tse_mac_transmit_endofpacket),
      .tse_mac_transmit_error         (tse_mac_transmit_error),
      .tse_mac_transmit_ready         (tse_mac_transmit_ready),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa),
      .tse_mac_transmit_startofpacket (tse_mac_transmit_startofpacket),
      .tse_mac_transmit_valid         (tse_mac_transmit_valid)
    );

  tse_mac_receive_arbitrator the_tse_mac_receive
    (
      .clk                           (pll_sys_clk),
      .reset_n                       (pll_sys_clk_reset_n),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_ready         (tse_mac_receive_ready),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  tse_mac the_tse_mac
    (
      .address      (tse_mac_control_port_address),
      .clk          (pll_sys_clk),
      .ff_rx_clk    (pll_sys_clk),
      .ff_rx_data   (tse_mac_receive_data),
      .ff_rx_dval   (tse_mac_receive_valid),
      .ff_rx_eop    (tse_mac_receive_endofpacket),
      .ff_rx_mod    (tse_mac_receive_empty),
      .ff_rx_rdy    (tse_mac_receive_ready),
      .ff_rx_sop    (tse_mac_receive_startofpacket),
      .ff_tx_clk    (pll_sys_clk),
      .ff_tx_data   (tse_mac_transmit_data),
      .ff_tx_eop    (tse_mac_transmit_endofpacket),
      .ff_tx_err    (tse_mac_transmit_error),
      .ff_tx_mod    (tse_mac_transmit_empty),
      .ff_tx_rdy    (tse_mac_transmit_ready),
      .ff_tx_sop    (tse_mac_transmit_startofpacket),
      .ff_tx_wren   (tse_mac_transmit_valid),
      .led_an       (led_an_from_the_tse_mac),
      .led_char_err (led_char_err_from_the_tse_mac),
      .led_col      (led_col_from_the_tse_mac),
      .led_crs      (led_crs_from_the_tse_mac),
      .led_disp_err (led_disp_err_from_the_tse_mac),
      .led_link     (led_link_from_the_tse_mac),
      .mdc          (mdc_from_the_tse_mac),
      .mdio_in      (mdio_in_to_the_tse_mac),
      .mdio_oen     (mdio_oen_from_the_tse_mac),
      .mdio_out     (mdio_out_from_the_tse_mac),
      .read         (tse_mac_control_port_read),
      .readdata     (tse_mac_control_port_readdata),
      .ref_clk      (ref_clk_to_the_tse_mac),
      .reset        (tse_mac_control_port_reset),
      .rx_err       (tse_mac_receive_error),
      .rxp          (rxp_to_the_tse_mac),
      .txp          (txp_from_the_tse_mac),
      .waitrequest  (tse_mac_control_port_waitrequest),
      .write        (tse_mac_control_port_write),
      .writedata    (tse_mac_control_port_writedata)
    );

  vol_recording_done_pio_s1_arbitrator the_vol_recording_done_pio_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_vol_recording_done_pio_s1                         (cpu_data_master_granted_vol_recording_done_pio_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_vol_recording_done_pio_s1               (cpu_data_master_qualified_request_vol_recording_done_pio_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_vol_recording_done_pio_s1                 (cpu_data_master_read_data_valid_vol_recording_done_pio_s1),
      .cpu_data_master_requests_vol_recording_done_pio_s1                        (cpu_data_master_requests_vol_recording_done_pio_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .d1_vol_recording_done_pio_s1_end_xfer                                     (d1_vol_recording_done_pio_s1_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .vol_recording_done_pio_s1_address                                         (vol_recording_done_pio_s1_address),
      .vol_recording_done_pio_s1_readdata                                        (vol_recording_done_pio_s1_readdata),
      .vol_recording_done_pio_s1_readdata_from_sa                                (vol_recording_done_pio_s1_readdata_from_sa),
      .vol_recording_done_pio_s1_reset_n                                         (vol_recording_done_pio_s1_reset_n)
    );

  vol_recording_done_pio the_vol_recording_done_pio
    (
      .address  (vol_recording_done_pio_s1_address),
      .clk      (pll_sys_clk),
      .in_port  (in_port_to_the_vol_recording_done_pio),
      .readdata (vol_recording_done_pio_s1_readdata),
      .reset_n  (vol_recording_done_pio_s1_reset_n)
    );

  vol_transfer_done_pio_s1_arbitrator the_vol_transfer_done_pio_s1
    (
      .clk                                                                       (pll_sys_clk),
      .cpu_data_master_address_to_slave                                          (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_vol_transfer_done_pio_s1                          (cpu_data_master_granted_vol_transfer_done_pio_s1),
      .cpu_data_master_latency_counter                                           (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_vol_transfer_done_pio_s1                (cpu_data_master_qualified_request_vol_transfer_done_pio_s1),
      .cpu_data_master_read                                                      (cpu_data_master_read),
      .cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register (cpu_data_master_read_data_valid_clock_crossing_ddr2_cpu_s1_shift_register),
      .cpu_data_master_read_data_valid_vol_transfer_done_pio_s1                  (cpu_data_master_read_data_valid_vol_transfer_done_pio_s1),
      .cpu_data_master_requests_vol_transfer_done_pio_s1                         (cpu_data_master_requests_vol_transfer_done_pio_s1),
      .cpu_data_master_write                                                     (cpu_data_master_write),
      .cpu_data_master_writedata                                                 (cpu_data_master_writedata),
      .d1_vol_transfer_done_pio_s1_end_xfer                                      (d1_vol_transfer_done_pio_s1_end_xfer),
      .reset_n                                                                   (pll_sys_clk_reset_n),
      .vol_transfer_done_pio_s1_address                                          (vol_transfer_done_pio_s1_address),
      .vol_transfer_done_pio_s1_chipselect                                       (vol_transfer_done_pio_s1_chipselect),
      .vol_transfer_done_pio_s1_readdata                                         (vol_transfer_done_pio_s1_readdata),
      .vol_transfer_done_pio_s1_readdata_from_sa                                 (vol_transfer_done_pio_s1_readdata_from_sa),
      .vol_transfer_done_pio_s1_reset_n                                          (vol_transfer_done_pio_s1_reset_n),
      .vol_transfer_done_pio_s1_write_n                                          (vol_transfer_done_pio_s1_write_n),
      .vol_transfer_done_pio_s1_writedata                                        (vol_transfer_done_pio_s1_writedata)
    );

  vol_transfer_done_pio the_vol_transfer_done_pio
    (
      .address    (vol_transfer_done_pio_s1_address),
      .chipselect (vol_transfer_done_pio_s1_chipselect),
      .clk        (pll_sys_clk),
      .out_port   (out_port_from_the_vol_transfer_done_pio),
      .readdata   (vol_transfer_done_pio_s1_readdata),
      .reset_n    (vol_transfer_done_pio_s1_reset_n),
      .write_n    (vol_transfer_done_pio_s1_write_n),
      .writedata  (vol_transfer_done_pio_s1_writedata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  SS_OCT_SOPC_reset_ddr2_phy_clk_out_domain_synch_module SS_OCT_SOPC_reset_ddr2_phy_clk_out_domain_synch
    (
      .clk      (ddr2_phy_clk_out),
      .data_in  (1'b1),
      .data_out (ddr2_phy_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  SS_OCT_SOPC_reset_pll_sys_clk_domain_synch_module SS_OCT_SOPC_reset_pll_sys_clk_domain_synch
    (
      .clk      (pll_sys_clk),
      .data_in  (1'b1),
      .data_out (pll_sys_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //SS_OCT_SOPC_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign SS_OCT_SOPC_clock_0_out_endofpacket = 0;

  //clock_crossing_master_ddr2_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign clock_crossing_master_ddr2_m1_endofpacket = 0;

  //pipeline_bridge_ddr2_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pipeline_bridge_ddr2_m1_endofpacket = 0;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane0_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 24: 0] rdaddress;
  input            rdclken;
  input   [ 24: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [33554431: 0];
  wire    [  7: 0] q;
  reg     [ 24: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 25,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane1_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 24: 0] rdaddress;
  input            rdclken;
  input   [ 24: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [33554431: 0];
  wire    [  7: 0] q;
  reg     [ 24: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 25,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash (
                   // inputs:
                    address,
                    read_n,
                    select_n,
                    write_n,

                   // outputs:
                    data
                 )
;

  inout   [ 15: 0] data;
  input   [ 24: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_flash_lane0, which is an e_ram
  ext_flash_lane0_module ext_flash_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_flash_lane1, which is an e_ram
  ext_flash_lane1_module ext_flash_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "c:/altera/91/quartus/eda/sim_lib/altera_mf.v"
`include "c:/altera/91/quartus/eda/sim_lib/220model.v"
`include "c:/altera/91/quartus/eda/sim_lib/sgate.v"
`include "Avalon_MM-Master_Templates/custom_master.v"
`include "Avalon_MM-Master_Templates/burst_write_master.v"
`include "Avalon_MM-Master_Templates/burst_read_master.v"
`include "Avalon_MM-Master_Templates/write_master.v"
`include "Avalon_MM-Master_Templates/latency_aware_read_master.v"
`include "master_write.v"
`include "master_read.v"
`include "C:/altera/91/quartus/eda/sim_lib/stratixiigx_hssi_atoms.v"
`include "C:/altera/91/quartus/eda/sim_lib/stratixiv_hssi_atoms.v"
`include "tse_mac.vo"
`include "tse_mac_loopback.v"
`include "descriptor_memory.v"
`include "pll.v"
`include "altpllpll.v"
`include "sysid.v"
`include "vol_transfer_done_pio.v"
`include "high_res_timer.v"
`include "sys_timer.v"
`include "jtag_uart.v"
`include "sgdma_rx.v"
`include "onchip_memory.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_oci_test_bench.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "vol_recording_done_pio.v"
`include "pipeline_bridge_ddr2.v"
`include "sgdma_tx.v"
`include "packet_memory.v"
`include "clock_crossing_ddr2_cpu.v"
`include "clock_crossing_master_ddr2.v"
`include "SS_OCT_SOPC_clock_0.v"
`include "SS_OCT_SOPC_burst_0.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire             SS_OCT_SOPC_burst_0_downstream_debugaccess;
  wire    [ 29: 0] SS_OCT_SOPC_burst_0_downstream_nativeaddress;
  wire             SS_OCT_SOPC_clock_0_in_endofpacket_from_sa;
  wire             SS_OCT_SOPC_clock_0_out_endofpacket;
  wire             aux_scan_clk_from_the_ddr2;
  wire             aux_scan_clk_reset_n_from_the_ddr2;
  wire             clk;
  reg              clk_50;
  wire             clock_crossing_ddr2_cpu_s1_endofpacket_from_sa;
  wire             clock_crossing_master_ddr2_m1_endofpacket;
  wire    [ 24: 0] clock_crossing_master_ddr2_m1_nativeaddress;
  wire             clock_crossing_master_ddr2_s1_endofpacket_from_sa;
  wire             control_done_from_the_master_read;
  wire             control_done_from_the_master_write;
  wire             control_early_done_from_the_master_read;
  wire             control_fixed_location_to_the_master_read;
  wire             control_fixed_location_to_the_master_write;
  wire             control_go_to_the_master_read;
  wire             control_go_to_the_master_write;
  wire    [ 29: 0] control_read_base_to_the_master_read;
  wire    [ 29: 0] control_read_length_to_the_master_read;
  wire    [ 29: 0] control_write_base_to_the_master_write;
  wire    [ 29: 0] control_write_length_to_the_master_write;
  wire             ddr2_aux_full_rate_clk_out;
  wire             ddr2_aux_half_rate_clk_out;
  wire             ddr2_phy_clk_out;
  wire             dll_reference_clk_from_the_ddr2;
  wire    [  5: 0] dqs_delay_ctrl_export_from_the_ddr2;
  wire    [ 25: 0] flash_tristate_bridge_address;
  wire    [ 15: 0] flash_tristate_bridge_data;
  wire             flash_tristate_bridge_readn;
  wire             flash_tristate_bridge_writen;
  wire             global_reset_n_to_the_ddr2;
  wire             in_port_to_the_vol_recording_done_pio;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             led_an_from_the_tse_mac;
  wire             led_char_err_from_the_tse_mac;
  wire             led_col_from_the_tse_mac;
  wire             led_crs_from_the_tse_mac;
  wire             led_disp_err_from_the_tse_mac;
  wire             led_link_from_the_tse_mac;
  wire             local_init_done_from_the_ddr2;
  wire             local_refresh_ack_from_the_ddr2;
  wire             local_wdata_req_from_the_ddr2;
  wire             mdc_from_the_tse_mac;
  wire             mdio_in_to_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 13: 0] mem_addr_from_the_ddr2;
  wire    [  2: 0] mem_ba_from_the_ddr2;
  wire             mem_cas_n_from_the_ddr2;
  wire             mem_cke_from_the_ddr2;
  wire    [  1: 0] mem_clk_n_to_and_from_the_ddr2;
  wire    [  1: 0] mem_clk_to_and_from_the_ddr2;
  wire             mem_cs_n_from_the_ddr2;
  wire    [  7: 0] mem_dm_from_the_ddr2;
  wire    [ 63: 0] mem_dq_to_and_from_the_ddr2;
  wire    [  7: 0] mem_dqs_to_and_from_the_ddr2;
  wire    [  7: 0] mem_dqsn_to_and_from_the_ddr2;
  wire             mem_odt_from_the_ddr2;
  wire             mem_ras_n_from_the_ddr2;
  wire             mem_we_n_from_the_ddr2;
  wire    [ 13: 0] oct_ctl_rs_value_to_the_ddr2;
  wire    [ 13: 0] oct_ctl_rt_value_to_the_ddr2;
  wire             out_port_from_the_vol_transfer_done_pio;
  wire             pipeline_bridge_ddr2_m1_debugaccess;
  wire             pipeline_bridge_ddr2_m1_endofpacket;
  wire             pll_sys_clk;
  wire             ref_clk_to_the_tse_mac;
  reg              reset_n;
  wire             reset_phy_clk_n_from_the_ddr2;
  wire             rxp_to_the_tse_mac;
  wire             select_n_to_the_ext_flash;
  wire             txp_from_the_tse_mac;
  wire             user_buffer_full_from_the_master_write;
  wire    [255: 0] user_buffer_input_data_to_the_master_write;
  wire    [255: 0] user_buffer_output_data_from_the_master_read;
  wire             user_data_available_from_the_master_read;
  wire             user_read_buffer_to_the_master_read;
  wire             user_write_buffer_to_the_master_write;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  SS_OCT_SOPC DUT
    (
      .aux_scan_clk_from_the_ddr2                   (aux_scan_clk_from_the_ddr2),
      .aux_scan_clk_reset_n_from_the_ddr2           (aux_scan_clk_reset_n_from_the_ddr2),
      .clk_50                                       (clk_50),
      .control_done_from_the_master_read            (control_done_from_the_master_read),
      .control_done_from_the_master_write           (control_done_from_the_master_write),
      .control_early_done_from_the_master_read      (control_early_done_from_the_master_read),
      .control_fixed_location_to_the_master_read    (control_fixed_location_to_the_master_read),
      .control_fixed_location_to_the_master_write   (control_fixed_location_to_the_master_write),
      .control_go_to_the_master_read                (control_go_to_the_master_read),
      .control_go_to_the_master_write               (control_go_to_the_master_write),
      .control_read_base_to_the_master_read         (control_read_base_to_the_master_read),
      .control_read_length_to_the_master_read       (control_read_length_to_the_master_read),
      .control_write_base_to_the_master_write       (control_write_base_to_the_master_write),
      .control_write_length_to_the_master_write     (control_write_length_to_the_master_write),
      .ddr2_aux_full_rate_clk_out                   (ddr2_aux_full_rate_clk_out),
      .ddr2_aux_half_rate_clk_out                   (ddr2_aux_half_rate_clk_out),
      .ddr2_phy_clk_out                             (ddr2_phy_clk_out),
      .dll_reference_clk_from_the_ddr2              (dll_reference_clk_from_the_ddr2),
      .dqs_delay_ctrl_export_from_the_ddr2          (dqs_delay_ctrl_export_from_the_ddr2),
      .flash_tristate_bridge_address                (flash_tristate_bridge_address),
      .flash_tristate_bridge_data                   (flash_tristate_bridge_data),
      .flash_tristate_bridge_readn                  (flash_tristate_bridge_readn),
      .flash_tristate_bridge_writen                 (flash_tristate_bridge_writen),
      .global_reset_n_to_the_ddr2                   (global_reset_n_to_the_ddr2),
      .in_port_to_the_vol_recording_done_pio        (in_port_to_the_vol_recording_done_pio),
      .led_an_from_the_tse_mac                      (led_an_from_the_tse_mac),
      .led_char_err_from_the_tse_mac                (led_char_err_from_the_tse_mac),
      .led_col_from_the_tse_mac                     (led_col_from_the_tse_mac),
      .led_crs_from_the_tse_mac                     (led_crs_from_the_tse_mac),
      .led_disp_err_from_the_tse_mac                (led_disp_err_from_the_tse_mac),
      .led_link_from_the_tse_mac                    (led_link_from_the_tse_mac),
      .local_init_done_from_the_ddr2                (local_init_done_from_the_ddr2),
      .local_refresh_ack_from_the_ddr2              (local_refresh_ack_from_the_ddr2),
      .local_wdata_req_from_the_ddr2                (local_wdata_req_from_the_ddr2),
      .mdc_from_the_tse_mac                         (mdc_from_the_tse_mac),
      .mdio_in_to_the_tse_mac                       (mdio_in_to_the_tse_mac),
      .mdio_oen_from_the_tse_mac                    (mdio_oen_from_the_tse_mac),
      .mdio_out_from_the_tse_mac                    (mdio_out_from_the_tse_mac),
      .mem_addr_from_the_ddr2                       (mem_addr_from_the_ddr2),
      .mem_ba_from_the_ddr2                         (mem_ba_from_the_ddr2),
      .mem_cas_n_from_the_ddr2                      (mem_cas_n_from_the_ddr2),
      .mem_cke_from_the_ddr2                        (mem_cke_from_the_ddr2),
      .mem_clk_n_to_and_from_the_ddr2               (mem_clk_n_to_and_from_the_ddr2),
      .mem_clk_to_and_from_the_ddr2                 (mem_clk_to_and_from_the_ddr2),
      .mem_cs_n_from_the_ddr2                       (mem_cs_n_from_the_ddr2),
      .mem_dm_from_the_ddr2                         (mem_dm_from_the_ddr2),
      .mem_dq_to_and_from_the_ddr2                  (mem_dq_to_and_from_the_ddr2),
      .mem_dqs_to_and_from_the_ddr2                 (mem_dqs_to_and_from_the_ddr2),
      .mem_dqsn_to_and_from_the_ddr2                (mem_dqsn_to_and_from_the_ddr2),
      .mem_odt_from_the_ddr2                        (mem_odt_from_the_ddr2),
      .mem_ras_n_from_the_ddr2                      (mem_ras_n_from_the_ddr2),
      .mem_we_n_from_the_ddr2                       (mem_we_n_from_the_ddr2),
      .oct_ctl_rs_value_to_the_ddr2                 (oct_ctl_rs_value_to_the_ddr2),
      .oct_ctl_rt_value_to_the_ddr2                 (oct_ctl_rt_value_to_the_ddr2),
      .out_port_from_the_vol_transfer_done_pio      (out_port_from_the_vol_transfer_done_pio),
      .pll_sys_clk                                  (pll_sys_clk),
      .ref_clk_to_the_tse_mac                       (ref_clk_to_the_tse_mac),
      .reset_n                                      (reset_n),
      .reset_phy_clk_n_from_the_ddr2                (reset_phy_clk_n_from_the_ddr2),
      .rxp_to_the_tse_mac                           (rxp_to_the_tse_mac),
      .select_n_to_the_ext_flash                    (select_n_to_the_ext_flash),
      .txp_from_the_tse_mac                         (txp_from_the_tse_mac),
      .user_buffer_full_from_the_master_write       (user_buffer_full_from_the_master_write),
      .user_buffer_input_data_to_the_master_write   (user_buffer_input_data_to_the_master_write),
      .user_buffer_output_data_from_the_master_read (user_buffer_output_data_from_the_master_read),
      .user_data_available_from_the_master_read     (user_data_available_from_the_master_read),
      .user_read_buffer_to_the_master_read          (user_read_buffer_to_the_master_read),
      .user_write_buffer_to_the_master_write        (user_write_buffer_to_the_master_write)
    );

  ext_flash the_ext_flash
    (
      .address  (flash_tristate_bridge_address[25 : 1]),
      .data     (flash_tristate_bridge_data),
      .read_n   (flash_tristate_bridge_readn),
      .select_n (select_n_to_the_ext_flash),
      .write_n  (flash_tristate_bridge_writen)
    );

  tse_mac_loopback the_tse_mac_loopback
    (
      .ref_clk (ref_clk_to_the_tse_mac),
      .rxp     (rxp_to_the_tse_mac),
      .txp     (txp_from_the_tse_mac)
    );

  initial
    clk_50 = 1'b0;
  always
    #10 clk_50 <= ~clk_50;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end

endmodule


//synthesis translate_on