��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t��v'gn�]o��in�m��+D(m.�B��/�����,��B	hI�ˋ������?�1J&�|WɆ&6�\]��%PM��t�&�m��'A>�:ET֤vKzL͊�q���B�s���e/W�������C��{����g³��ws�#�=ѧ�y�A���Lc�����Ǯҁ���Δ�'�1�����7 rG�q���(Ƥ�i�Q����`���?H�v�d��]oDO#���Jꘜ5�1��4�XUY�����N�Ae�#�����B�N�By3��<�]�!��	Ǹ�y85�;{��T֧�6��	���`y����ꢤ�Og�y�1a}�c��Et�Y�{'%s���䒼�W& s�����"X��[��Q[R�7�M�g����Y%T��BPe.��xu	�>��l%i�-��9��稕Y%T��BPe.��xu	�>��l%i�-̇i�d�?�Y%T��BPe.��xu	�>��l%i�-D�wP�/�wM�Ǿhm��@IE�U����S8�
T�F���u�܎����k/��m#�U��_D��.V&��B֥�(����5��ٌc�5��8����Bp}|��XH��9��p#�7ڜ¸<�X���(����5��ٌc�5��K�E�\��Y
iEE�G+�T�J��h�H�MPq6.�b9�����6�_��1�m��'A>/y,�Z���rS�b�8Z���'�e�����"�?;(��j67�=t�!��&r���q� N��p����IÙ=�Hʆ�In��t/p���xL��fl���=��fLR=t�!��&r���q� N��3�AŠ�zL͊�q��٘�27!�g?_��<'P��!jcCA�T�g�v����fQf��p�m~|��4FV�{E�JHn��z�'8^�#ٸ�U��֜��3Ԓ��������\6��.�E�]��c8?-+eN�s(^��^p��nk�Y�P	dU�1�1�����1#��Z�����XP�����'�e�����T�LJ�n��f�e��}�
�?�`<Y��sp+N�f�+�n`5�fK��0z�cUL�?m ��0���k��$a(􆿳���2����.��DP֞ �T�'Y���A�? ��p�]�!��	Ǹ�y85�����S��Cƃ
ᾆ�x�T�\ ��i3�|)sՀ�T:���V�Z7����6	зq8�Ј'���Xw�j�7��Po�Q�>°������R�wX��}�
�?����2jɸ4�r�@E�n`5�fK��0z�cULn�4Z_U���l�����"X��[��Q[R�7�����bpZ��	�`DÜk�K��h�d�٣��c�A�L'�"��/f~�\	��K(����`y����@����gG�������E3-	����#�6�3��rs�i�_n����B�Pcsù��Q��Y����2����..W���ۗ���WYHpYyI|*����]�!��	Ǹ�y85�����S��C\	��K(����`y���_���e��� X��V�+�3q�bx�#�;� L5ӥ����S�ۗ����f��DE3-	����o�?{/T{9��#.���G}�j�d�t%>^�ߦ��|R%��<��0n|�!h�b���t�m�+�L�w�s+�¤]�o"�s�8��cEp	���>P�2-i_q?�y��T֣[\5qJ�}���2�WaU�W�"c��ƃ
ᾆ�x�T�\ ��e>۵��>��?!6)X�TuHuJ����V�2�R;+�l����؊�.�����ӯIJ B���J��>���@]KZ	��\#�Z7����6	v{��lw	B�*
cR�'6���;8=�g��U-�eӢl*H0*%�W�%�K���ⓚ�����>Pcsù�NdE��Q���;mQ��b�c��=9�ߨ�,R�A�=��Byw?��|��ՕH;u�o��_�Rv�䩲$���dS@Ɵ�o{y����i�q,?5q��C"�M��5�:��\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�D�wP�/�wۏ�:��"�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^xjzӝ�������iPo�Q�>��aIO-�����&G!�`�(i3p�n���/�i4?$|�ڗ�\���qhF�fp�Z��	�`D�\��v� H���;mQ��8���/���}Dq�f������!�`�(i3p�n���/�i4?$|�ڗ�\���x�o"jU�Z��	�`D�\��v� H���;mQ��8���/���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��C"�M�4����(��5��
�c�{�#�I����~uZ鎬�������(����.��$�ʝ.�&J�!-B=�6f��Z:S����b�Bϱ�O�E�l`8x뛀���!���"��o_B�E�JQm��	�̷_��yC��S8�\�w�4�'�)�Բc��?!6)X���%A������D�ϲ]�6��2�S�i����T���!�`�(i3!�`�(i3!�`�(i3!�`�(i3��>��lJ���aٔ^?���S�T*��;1�˚�!��JlR����2jɸ���[=��u���������-��d�XS��_'���Xw�j�7��AԢ�a\�#P��W��������|Pcsù�u�ȭ�>�W��7(�bOI\�w[���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�a�}�$��W�6?���N��S��pP�Fc�����k��$�����k�A#�G=�Yկ����!�`�(i3!�`�(i3!�`�(i3!�`�(i3��͉��@��B���RWL~΄gO�3��|��[�侰j���