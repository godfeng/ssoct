��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:�� �c�=0N���6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,xh'�$k�w�D1���}����ň���x�w�Y��k��ı���$��������j��t�w )�1��kN<��;��� B]�pE���	x]̃Dj#^Da����M�ٲ��9ߪ�
�M��ļz����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��Sd,�ϱ����@N1�w�0XL��t:w�~�gm��+��9��kT!����Y�f��a�Z��V2 �Q[6�i��<&�̝n�U��Y�C���t�#K�{ʓ��d��?�A\���5���a["<7U�i�#6u�,Уd�^:$�$���?#�+jN�N�{M}@���x�h�v[�2)ݛk�}dXQ������K����{Z�/*0�(bѮƷ��,�&'��Y_�68m}C��Z1)fd�vĻ�E����F5���Xf/���Jm�WH)5�Z!{����
F�P?_�!B�]M"Aw��-��ׇӭ��!�`�(i3!�`�(i3u0��L<q�`�c&�r.�?cXE;�i~p��M��gCu(o?C�����5	�)kJ#��t�{ڼ�`a3� �x���f:3���/�ky3�����=��ׇӭ��!�`�(i3!�`�(i3*8�2�z�����b/?�8I.���^r�b(�c�?����4����o���������i���%��S��!����P�><1N��r'�)d
�u|�$�iah7��f2`�r��sȸ�"rR!�`�(i3!�`�(i3R����G�ތ_tO~��E@�͔��Ġ�L �*�2R�W�~�26��\K�y؄@�!�`�(i3!�`�(i3/��oi�#��+��:iR��Sp㨚��}��6�8�-Zy?X��?��W���;��B�lXK�y؄@�!�`�(i3!�`�(i3�Կ���pu&a�vU0��p�$;�n ��j�ּ���)`4Zp��/���ϲ���>h�c}����>I	���(��B�:����@���4W�-c8��"3���s��ׇӭ��!�`�(i3!�`�(i30R��=	�@����W��nl@O4茸z���q����R��C���CS�� ��!�`�(i3!�`�(i3�0�9&،EB����n��|1�b�YL��&\VI`,xJ�����g}����&�������!�`�(i3!�`�(i3�>=���#9����'*�J�.�����G����%�,b�_�Ќ��*��4.���Xt�.U���ͧ�uQ0�})�����,]�x	��gf���{�P�1|5я����j���ֵ��sȸ�"rR!�`�(i3!�`�(i3_|?k��\+X��Y��8�-Zy?X�!�ZN9���2�䦒ccnh?�!�`�(i3!�`�(i3��j0��x���jz�H�gf���~�c��"��&\VI`, �DO'�L!�`�(i3!�`�(i3����N���z�����6u=�{��ZMN��>�! ,��e�w�1V�N��:˽�_k[9��~��!�`�(i3!�`�(i3'�Z�8�'��ѯh��d�J�\���=��&\VI`,f���a�9e47�O��C��_���U�`�R�Z-��شУ�X��d�rW��y����Fz�!�`�(i3!�`�(i3q<m6p��*u�j}@�El����WtUr���dp�
�2 ��Q=ߎ�����,������ccnh?���&\VI`,�=JK�t�J%�r �14�X#�Mwn5�����z1�z�F���ϡe����W*�RYS�Kh�!�`�(i3!�`�(i3!�`�(i3�q��L�!?�d���&�u&a�v��� a�ik��Wʍ3�V�޷��i�mm	�>!�`�(i3!�`�(i3!�`�(i3�@��ÂbݩJ�\���=��&\VI`,门:<#B�����+C���~KM�gzu4��	�!�`�(i3!�`�(i3!�`�(i3�U��a��*��>i�!i�X!�!D��(J�f�)�s�%�hH�oe��C��c�S+d�J�Г��f�u�����!-��B<ԧ�[��+��sȸ�"rR!�`�(i3!�`�(i3p{���gM�k���lh�&ĵ�	ƹqE_���RQ�
�)T^�b�k�@����S��l��ׇӭ��!�`�(i3!�`�(i3J�Y,�~)�{lN}Q�b�o�m��}�؝�TVq�|`kK��I�t����ۀ ��m��5ѧ��Z>)E�d��Z�����d�*���Fz�!�`�(i3!�`�(i3������!���C�/�y���ܴ�WM�P[��j�$�*7I���y�L�=sȸ�"rR!�`�(i3!�`�(i3+���6>�2'5�sZw��Q����}2M�; ����������-N��]�1�l0�)�Myիnň��h����]ߺ�`@��h�h����M����CN�u!�`�(i3!�`�(i3!�`�(i3��_�����v�����������U��5�D�v�l�Ū�TD���wG",���˫�i�m|� ��>K�U��L��nc�^��ns)��E�$�S��Z(�j�!wS����G�N�����ڭ�[��
A�4ϦE�6����ѹ��6[��{ֱ@����G��Mr�J�Mۀ7���\� ��2Rn�k�*��� ^ȣ�2$6�sI4$2�¤}@|��d��\��'ٽ$Id`ȯ~���Uz���+ߜ)��ns)��E�$d??�A��?U��|�����X�4V�.�(A���C�/�yV<��ϚEP�@�z���c>�I ��bv.�]0�[X�b\g!"�a$��z�e&Y��WM�P[��=����Vq�|`kK��I�`\�L',�y�+(̇�0S&",f�e��sƲ����e:ɄP���'㦡���0�8*��#�N�J���}��R���j�y���i�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������ݧu7Y�M�+|�#��Byl}Vİ�8�d��N��Ԫ^��rL�t��^�:AԪ^��rL�g�j�m��}��w�G���RJ��p�99-#` ������b_]s��2��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcfe./��:�!9\��N5�w��J��Zo  �0WP�da����'Q�:��~�z7	9��sE���ye��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#�.�x^ok��u4�� L�ʿԪ^��rL�Nl�Dvg�	Ԫ^��rL�t��^�:AԪ^��rL�>���x�<Ԫ^��rL�%�7��Ŀ<Ԫ^��rL���7�C)"�Ԫ^��rL���	��D9�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcQ#�y�&(���B��|/~.)��3\�R�F*}�c}��uO�^VM,q���\��K[�J�#��9�ĒTC��0���^S�kC�"�Z<�
�#*t�uADa��?4j��a����2�˴L�t#[����p������*�۽�.�jI`� r��F'�J�|(�����	x]�V������g��Z~Y��]#�]E���4������D��a�,F�7&�����pN�Wu��w)�S���f��^@�~篟|�Q�M�u�c�.C�g�dџ�_�v%��O��J�O�� 0�^"R��#'5��i���~+�lX҉ys��3Tb�����?�����$��w���މ�r�O��C��0��QP路h�����G�/9��g��G��������!�zg�Z�$�����j{X� ���
� �AH��1�����Cn���ʯa9̷�
�Xg���e�JrtΣ|Y���%�����φ��~��➛����T8�{��3!Z�*_#a�/����i���7�`ѡz��9���vo���Q�g����#$^��j8HQ��X�t�q���ѧv;��gf����)F�Z�u6_���͌�<�vd�̪?�d���&��P�>�� ?[n�:#G����8
B�ɹ�`S´ c��(�U����	x]�<��O~��#?���/��di���� J���<���&}Xa���qd��.�wjX5D	1%���n����k�8���҆�|n����﨩R���i&��a��fx���$�U��"�>�q�ax�MU�٣�R�B;����4G�n�?�`7�K�|���g�3] ��Jkŏ��8%C��c�S+d��t4�f%N�XG���\�4�s�q�=Q��xY��݅ 0��|�~���nM�bb5�Sd,�ϱ�ϖe��!I�I�� n "<W55��XR
ئ�v�5ܗu��S&ϊHF>iDj(���ʇ��p��x+65�p����o L�"��\�4�s�q�=Q��x�)�����|�~��wU�����Sd,�ϱ�ϖe��!I�I�� n "<W55��XR
ئ�v�5ܗu��S&ϊHF>iDj(���ʇ��p��x+65�p����o L�"��\�4�s�q�=Q��x
�ԟ�d�F�D�Oo������o?�M��;]�;��
<�����&��*�_��l��f���<zT����H��6Ó�KF�vw�}\yȺ(��m��A� c��(�U����	x]�<���e�0�9�(��`ݓ��� +u��Ipc9�`s�S�͔�Rټ ��߷��\�4�sR���i1�8Y�&�\���p�h�%ģ�l�$9Ř��W(�1���z���D)���pH�P�SyH�O(ٛRF�",�uJEA�����X�(c��k�8���҆�|n���u� �(�eg>��rvp�){�~A �ѕ�����aWfL1�;4�zu%�1<�$z��n��kF-�F敪29k~��e&~�:u��w)�S��X3���7��Mv�9����Dtr/���zbl�џ�_�v%��X�'b�mh}����N�@N�����N���6[�'�&�' �>�u��8�F�D%� ,R�w]�y�ljrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;�m�\��qi��p�7���I�4��ʆ	��i��p�7��Z鎬����~x���i���;t˩�e�J�4>��1lD�J8���=Udq��D��tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"~����d!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������N{a�9Ow�Y��k��ı���$��������j��t�w )�1��k�+(��<UC;6aJVlO/������V��r:O!�`�(i3=]A��O�T%��^[~p��M��gCu(o?C"�,�>E����\�v�T?�7G|`��#Զ.���@����!�`�(i3�b9���:&�>��s�4zG&/���o���������i�%Ah�%4
>��XP���^�Bmw�D'�H��H�8�-Zy?X�!�`�(i3JHn��z�_c)���8Л�L���P��}��6�8�-Zy?X�%Ah�%4
>��XP����@aw��r�],Aبs�E���-{o-�<<��89X�������B"�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD*�\�)M�rO�N�U�#�&0J7w� K8�&+1@�D+`uώ�:�O,�у�i��؞�x z�Jm]A�/�����%>%���P&c"����Q=ߎ�����,����7�ܥ��2�� z���@��xR�"�,�>E��4];ˍH�!�`�(i3���14�:v~E�)d,^<���cO�1�9��`�ox!�Q�W���`~�ߪ �)	�8Vt%v�
�9�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��J� �Y��0�4�+��V�-��	�G[���#�4���Wj�6���}2M�; ?9Pjp���Z\�+)epl0��F��j0�T��:�wH�HͶVq�|`kK��I����+�J��U<o^.K�}�sђN�1�c��N�w�Q^�MY:��]n��JHn��z�C�$��؍��R��j�.(Wx*�_F�k-�!�`�(i3��|g�Y�'���Xw�������펎��{5N�By3��<�]�!����M[��ǢK�h-L���H�B���5�¬����"�����E����F��j��\w��0]vwdI���<�_�r�)�s�ި�(@X~�H:#�<���Е�(�
t�ژq���U�[��N�霬�^����Ú���Z鎬�����	�7 �#�����g�0ˋ��I��w��,>����C��(R\֎u�3�i��7G#+��\w��0](@X~�H:�+�w>����(�
t��Y�{'%s=ͱu���D�v�l�Ū�TD��������B���xBP��_c7�v�ԯ��Q[R�7a�s�9���)Հ�^2��b��|2�����i�M��cg�P�TD���rs�i���`�M�	=̞��>�B^`ٌ��x�[5��Z�8���/��?uF�Cg4�Y�J�Yl���#�]�!���D��L#�����/��]o��in�m��+�<4��ˌ�ň��h��j�V��v�����>���C�Y�)�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�L~΄gO�3��|��[��"�Q:�{�1k�ZV"���:��#tC������s�Q�_;�"l���Bp"	���@����gGy'q�;�����Zv���;�b9����`�Z�kU�u<^�T+�B-�D ���3�Һ��7U��sb!��u�-��>lf+�S���c,��\�v����,Df���	\FX���CUM��n`5�fK��0z�cULd�g>57<��ʹ�q鳏G������W�\��`y����@����gG=%� g�Vv�5)��Z^7s�9���o>��l%i�-5�e`��9�\1^O�cɴɫݜ�Z鎬������_�,�[/�cWM��@EZ������Q]� _ό���.�}�
�?��Pۢ����!�`�(i3�d�٣���N N�S�\�#$�ÙA�,�&Ѷ��зq8�Ј'���Xw���RY��EOJ�uxm�v�����;�L���9�f����؟�r�1G}�����g��U-�e��,G�#�Y�{'%s=ͱu���˝Sz��E�4.@�7��y%%��`y����@����gG_�l����i�N�.�69�<���v��������,D(q!�_�{&Ҽ�q��]�!��RY���ت�`�������H9��p#�7�Q,[��;!���v�Z��	h��4���b��M!�)HnvKr�3�͉=�?��3��J��R���=�?��3�w�kZ"�jX�qp�c� �`p�~(�M#�<���Џۢ	:j���1�, �!�)HnvKr�3�͉m�a�gPM�I����~u}���yb��H9��E	E��BLV�v6�#�����i7N�_�wDo�h�'�t�Z�f�}��+��\��5��,bXh��d���!i(@X~�H:L�����l������Ho��'�\�n`��!��BBaYz+�Z����~R���1��� ����P�7� v{��lw	N�]|-�ǳ��&Ҝ���,�ǰ	M,��rERj�V��v�Z� >�
�,�&�X�<x!�g<~�i}VCk�HtY�S
�I���R�U��)���Pa�L���쥗>�Ϳ�F�� J�ʯ�7I���VjԿvU!�`�(i3�3FV�J�3פ����t��}pshI��Tޅiy:Vy�a���$�Qu�|�E �jǳ<��C�
�E����F�5F:	��ֱ�q���Q��^��N�m�[�N!�`�(i3�d�٣��c�A�L'��~�2�?�B���N�gl��ܬa(􆿳����^���~�26��\2|Oo�{b�!�`�(i3�rA���oq��WX ��b�FP&���Y�l,��\ُlT5�i3<�f�D.`�Z���N}�m��{�Yg3J���e둼�;зq8�Ј�)V4�$�!�g��U-�e��,H/�� ��b�FP&ӝ�9��,y�
j�m�f70���x�]�V��/��A���U����I��N}�m��{����g�	׭C9*�¢�������r�Sy�n�yLjn�=m�"�2N��n�[�hŽ>톛z~$���"�,�>E���"5� �S��s��?�2N��n�[�hŽ>�h*�t�8�N"�,�>E���"5� �St-p���|ȧ2N��n�43bXD�O�$&�<���c��+)3��#�ڊ<?@o����δ��q��(&�L��'ž1�|��P�:k& ��-����\���F�`y,�[��$�w<���x�����*ȑs��-�����y��j��k���J�4�y��Nկ����}Dq�f���Q��}	��oo�@L=�ω.t��U~܎VV��.��J���&_��=]�RCJ�����@�ĵm�ݚ�Н��]��/ݐ������YF%�"�Z1��2�A�dv�:5A��p�)��S�2�oo�@L=�f��0��o��!'�1tSjv��/��@����*��Sx�m���n�>�<���x����:5A��p<�6�Q=�����ټu��.t�5�M�1�>�scX{�X!,�wbk�$����$�Ӗ��Y�l,�~ov7#}!�`�(i3���gRI/��K�p�9"ʝ���ԃ`!�`�(i31���~���y��lDR���1w�������c�I���8��1	/�!�`�(i3M���COp[U;� �M�[����i�u���U�Uܲy>!i��{�.D��Ea�7㑠h(W�y]�2/U �t��]�w9"xO��S!�`�(i3�8�ܩ�ò�]�B#	��?D�8��9��n�7�Y���X�q^օ?D^��!�`�(i3NY�U���Ȓ�m���B�A��o>U���b�|/B�/?�+t�<Ǿ���������~����p!��
`ϙb9�O��F�����~}>�O���(
�T�r�5�9�O��F�־^N��ܱ�{1?�a����h˕��3��a�-$�x���=��:5A��p$f��_Ub�F�S�1 ����F��O�t�{#	�x�O�M:R	���hIf��{_8�Y��M��)=໺(ӈ���]!MuV�	���̰�!w���B}�#QSU:�����|e"���x8�!�`�(i3%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩη�X��n�;��0C��;g��&�����6,��$e�<O���,9x{^4��*m!�`�(i3�]�.�,���9z���@�oS��ܠ�a�,��
�T�r�5�����l���\�A'YE��"� _̸ ���]�0��Olz!�bf���,�����Qf��� :��
&T��'���d1tSjv�!�`�(i3q�ޖ�v
>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ���Q[�lm�>&S�XQ�������x{^4��*m!�`�(i3;�jmT�#����n,��>]��e������Y��7����!�`�(i3!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3!�`�(i3a�/�	5�{1?�a�/}�׏)#uE9�+��!�`�(i3;�jmT�#Ό���;���P*e�{�W!�`�(i3!�`�(i3� ͷ�	�%�s����V���a�٨���bN�F�!�`�(i3!�`�(i3F�Q��^Wp��9B����U���uE9�+��!�`�(i3!�`�(i3:�HCaIMl*h~U�?u��l(E$3Eur��9�C!�`�(i3!�`�(i31���~!�`�(i3�/��@����*��Sx֐�M�4m��?�N����!�`�(i3!�`�(i3:�HCaIMl*h~U�?u��!���c�A�L'M�M˫ɒ�1��!���1Uk���D24N<I8����\.W��v�9��!�`�(i3���%>�rGO�D mWN!�`�(i3!�`�(i3ѠZ��<���l>��~�
�aLS����>�)֚�I��&k�F� w^��t����v�q���r����!�`�(i3����Q���~���c�6�fST��*b.[P��=���f.K!�`�(i3�H�����8�ܩ�òo�����=������&G!�`�(i3!�`�(i3�<�W����6	D�NQ�4Ư�ƧE�f�s�#>������!�`�(i3fĉ>99��A0ok��!�`�(i3fĉ>99��R�Q���~��p����!�`�(i3��w�w:�!�`�(i3!�`�(i3a�/�	5�{1?�a�/}�׏)#uE9�+��!�`�(i35�����}Yms��/�u���4���O�>�k}�r�,0=]^	�&��|�B�����Yk��!�`�(i3�,:��#��@��xR��_���1tSjv�!�`�(i3!�`�(i3���W��Ȑ��dȠ�$h<���WㆴYƨ@0�$!�`�(i3�?�W/)G~�`cC�4��.��cZ������N��}Dq�f�!�`�(i3�2��}��E2�DZ���  ����'c��ʿk�M�|9��zD!�`�(i3՝� s�#���k$ !�`�(i3.��J�޺��:p~	E�<l��uE9�+��!�`�(i3�2��}��E2�DZ���  ����'Z鎬�������(���/%Z�ڄ^1[]�]mu�5v��v�K��������ȓ=�^݊��}Dq�f�!�`�(i3HN��R��bP�63Z�t!�`�(i3;�jmT�#�B�%3�Y]�|�$�&�U��f�!�`�(i3!�`�(i3�r'Z1p8j����I~��;��7=��9w�ƖF���m¡!�`�(i3���%>�rGO�D mWN!�`�(i3fĉ>99��R�Q���~��p����!�`�(i3$f��_Ub�F�S�1 �!�`�(i3�(R\֎u�eK�	�$V�n��뾦�!�`�(i3HN��R��bP�63Z�t՝� s�#���k$ ���y��lD�ה3UF�׏23����.L���M���i��C@!�`�(i3��;��L���W��7=��J����;4�zu%��5)��Z^�'����u��r��!�`�(i3�%t̓�@��5)��Z^'�^�����ݚ�Н��wӨj]h�O�M:R	���hIf�套�qD0�5`�JBu'!�`�(i3�����!�`�(i3ݑ���&�d>&S�XQ�<F�ڴdƍ2���l�!�`�(i3w�����A��N�.�E�g����������y�e��0�U��JeR�&�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp'{w#/ B<�6�Q=��ԩf��Z!��
`ϙb����l��
*kB��`x�W��7=#o�]�ʄ�;4�zu%��5)��Z^<���H ��;՟��1�, �[���*1tSjv�!�`�(i3���x8�!�`�(i3n��뾦�!�`�(i3���̰�!w���B}�#QSU:�����|e"�wӨj]h�O�M:R	���hIf��{_8�Y��M��)=໺(ӈ���]!MuV�	!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M;�Ղ���-,9��-m��-�$��S&ϊ*7�xs��^	�[0
��o#��|Zb?�����&*; i�V�JD�IX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>���9�.J?�(z�)�#�xjzӝ���w3��׍�&�U��f����1� �.�
�ɺK� |�>��̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^oв%u�K�>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ���-����!�`�(i3 �bVfj��h�c,.J�AԢ�a\�%o�P��(� ��0� 1tSjv�!�`�(i3?�����&*����@z\��}Dq�f��	��x��ݚ�Н�џ�3~�l"+�B-�DT����?.�s�j��0>������fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹��x/�Nn��&v��;}it�d��"�A�S[W��ցDG��X�"z$x�_~�@Q��mU�ߏ�˯�h"E&��� �n9�O�k�*$%M�֞NP���G��U��)���Y;e�iK-pm!9�>�k\������`�5�i�+�؟6u�0���$�Qu�|�E �jc|��U�	�I]����2N��n�ܖ �&��T��opU�ތ�K�J���N}�m��{��F_��R�%�&`�������o0H1��M.��jJ3�9�C�s�4�2N��n��bcb�q�\ꉂ��dC�&T�F�9Ặ��Ϊ�Q� ~��d�G}%����3f����;����*���ShT������qD��=a�^7�1tSjv��A�Z������**,n����"� ���c�d�1��Z����<�>�y&	�eu�o������?�&=q��m�31���,��8�-Zy?X�{ݮƻ�@@o�'�P�o�BH�n?a�1#܆<ȶ}������9�O��F�־^N��ܱ��*����׭����WI��0�4�"����-2w ϣ酋x�Ifl,[�跱�:�윯}Dq�f���m�5h1��s��Xuz���_�o��p{{�;ͥ�H�RtV�^�: -Cx䪌Y�6{W�(�]}Ϳ�#��̢i��;�C���E��&\VI`,�=JK�t�.��$�'�ͬ���~,�H�͛�՝� s�#���k$ H������r��\E��6f��+�<.+6J!���%>�rGO�D mWNHN��R��bP�63Z�t����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l��	ͰZ����5)��Z^�d��-��!��KVט$�W��7=#o�]�ʄǸe�q�A�ވ��*I���b�Bϱ�}���yb���?\MP!� u��r��c�@�/��K�X���X�y?-O딈pᜯ}Dq�f�=q��m�31���,��8�-Zy?X��f�8
��u��r��!�`�(i3r{�"���.ޟ���T��=y����͘6��q����1ig!��v�9��!�`�(i3�JO�'�����n�@���^����!�`�(i3a3@��[/�-=�f��W|N�Y������f��`ȱ���}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}ĝ���;����*����nûdI0L$O�a��Q��\�"ߗtˍ���!�zbf}߂���ȍW�����I��.ŭR±���J�q��tV�*}�S�Ҙ��3�_��Պ-�ð'տ@x��y'��BS��F&ѐ��ŁG&y��9�nC��s+�d++~�S2�h�φ��<�6�V-T����N}�m��{����g�	׭C9*�¢������7k��/j�Ch��㉊���;���EWr�c�Em����<�u��s$y�<H�-��*N}�m��{�`{��U	�f70����W0i��^O��bvq�ֱ�q��WaU�/G5��d�C�U=��W�E<HӍ��`���oN}�m��{|�v������!���JHn��z��
�kˤ�:Fa�7�����PϾ��Xmt�=���3��a���!@�f")u��r���**������fg(VQ��v�?i�:!�`�(i3-���H�� �7~�	 �b~*��s��(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<�QtOn7�\!�`�(i3��y����u��Ƌ3�(R\֎u�eK�	�$V�eW���Z���I���!�x=�FZ|V��K�ѧ�4.���A��F��ݚ�Н�(*�O�q��=�����!�`�(i3���������6�f'A��x�x�]t�ݚ�Н�Z��JP�����>�Q��!���c�A�L'W»��`�{�L�de����G����vq����ۉG�e�&&�����/��3��}Dq�f��mJ�0�6�!�`�(i3����J�V!��d!�`�(i3��z�Yh�ü����&��2��M!�`�(i3����(L֡��|W�֨r������)c�S�l.|���!�`�(i3t�2E8^#*��*$2V ;��8�q<�v 8��o��+eQ�����)M��ݚ�Н��� л��x���u�&;��I�H�^&s�����*.!!�!�`�(i3�����i���@]
�a�(���B���Oo��[*��������:5A��p�0�9&،��F�z�8#��%L���rS�b�8Z�}���yb��CN�zB�!�`�(i3��t��k�b���N��B�4]������@}➛����Xw�e60���ǂ�e��sHb�����
�!�`�(i3���Q�| V�}zj>�c^g��G��'r=I4�!�`�(i3��yl���^�K�d{��8ѭ�B@s�tY� h�ҩ�!�`�(i3��N�T?w�\�ϕ��dW� g�[�܀Y�I��!�`�(i3���F��O��ݚ�Н��H����jF�ཕu��Va�ir�8�ܩ�ò�CFy��Q������&G!�`�(i3�� л��Vr�������ltY��1d��mw�x��F�;���!�`�(i3O���8z����( k��o�{��Ļ�*�@;��-b�uE9�+��!�`�(i3%�yLp�h�C��_U]����9�suE9�+��!�`�(i3Q7�.2B�*���B���{?��ބ!�`�(i3���y��lD�6[�O�?�f��!��u�M�ｂ g�!�`�(i3��z���>�-F�#@�����F�z�8#_k�B�a��� h�ҩ�!�`�(i3�H����}���yb��1P.��d���G����4Xf��GH�RtV�^!�`�(i3H�����?�@,��Vҙ2�f�������]!�`�(i3!�`�(i3��Ě�����}Dq�f�!�`�(i3��Ě�����}Dq�f�!�`�(i3�5ߧE4��!�`�(i3H������B2|X��̷_��yC��S8�͍u�	�g؝�b�Bϱ�}���yb��/�!U�*<=�*�$���i5{��s!�`�(i3�̢k������Y�l,��P5��"G� ����v��f��;2�5�p��`C��Y��H�RtV�^!�`�(i3}���yb��r)1;�Os�rs�i�}�O��L��_
�u��U.+"b4!�g��K�,>0���0��Jn��ݚ�Н��/��@��k=�E�ɟ_�ܾ7�'�� �����F�V�hU!e�Wm�r�ʆ�In��t[�(����W��F�z�8#�:5A��p
�:qEp'{w#/ B!�`�(i3��vq�|W�XX�<f�KV���a�;�Be�\R }��i��3�!�`�(i3H�����?�@,��V��\ �I3�|�$��N�u�48b�������}Dq�f�!�`�(i3}���yb��s��O*m]Z鎬�������(���Y�&�-��Oj�\Ʊ؀�o�P�}���yb���}��0�X��v�9��!�`�(i3M���CO�0 ��%O7�9�u�����
F��<�d��@�&�1���"�A��K��YF�"�؃l��J���֨�{�Y�!�`�(i3HN��R��F F�E̠!�`�(i3������I��~�Tz!�`�(i3a苯ܪ�\�k4|��1+�M�r�r���S���ݚ�Н�(*�O�qe��0�U������K!�`�(i3��4�CD5���}Dq�f��5ߧE4��mJ�0�6�$f��_Ub�y��D�nmX�Fr��j�@�f�smy�zԴ�	�����}~�.���
�y'��BS��-��%j��Ak|ņ�R��cÇ�ߐ�*��#v������ ��M'gag�bR�jZ��;yE�f*��$-�p�ny�(H`��Prm����6>Յ��ogg St�T�bCJ�L#��K!�#n��]mWᅫw�5�O�%E#P�$��Xo�<�OP���-8p~�b9����r*�^�	�?�9IU<6�N*;|�m�0�l��*Q� ���V/��w�i/��T`�-�	B(�	<^��.�Q�s	���0������v�#��s��^g�)�.�z���g6�^g�)�.�I�WO`���\o�LCd�w�[������v�ł8�cB����ʢ�����8&���Ie��  �Í�sr�>u�quA0�e��^�uJ#����+�^n=\f�5>��9��mǥ�|��S���R��%4��"S�#�vzR5�<��b+}y[i`YS����Q�޿�ߏ�˯�h"E&��� ��!�>����T�z�)tŸ3y������UTM�Xt���p�`ݬ1�N�D��泵l�QR� #�R�U�R��8~e�o1n ��F˷^����o�����?o�#��J�g[j�"2xM{�@c����'R�����z��_���mA��$}�O@���cB�8� ���'��������լX�����%������������9a[�-�����4�Z�Q�D����4q�.-�gg$�/bKCEɆ�SV"@]��2Ƅ�}�U+�~="�����:��ȓM�Me�����(�z9a�<�Vr���1�B��aU�1Tn�B
'�����tl�:�K*��gB���A�_A��N�Z�k^��0E�Hg������n/L�D��$������A{4}�u���_�A�|����R��%4��"S�?�����&*rB�WD�{͘6��q����1ig![ �#�|f;4�zu%��5)��Z^�d��-��!��KVט$�W��7=#o�]�ʄ�m�Թ���p�T��~��d�>���{#���J�������
��'1�Z�)QvZ�P�C|���дV�fL�V���_���{�6�C������n/��V8zA�o��<���� ��V��G��<��
��)����y�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�F�KD�Vr[/}>5��0+�_0c ۹1�)��ٵ����
�{�+q�R9���Ih��Z�)QvZ�P�C|����k��.���SxF��s���D���{�6�C������n/��V8zA�o��<���� ��V��G��<��
��)����y�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�F�KD�Vr[/}>5��0+�_0c ۹1�)��ٵ����
��Viņ�9���Ih��Z�)QvZ�P�C|����k��.���SxF��s���D���{�6�C������n/��V8zA�o��<���� ��V��G��<��
��)����y�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�F�KD�Vr[/}>5��0$r�t�}i$�)�vx�9��m1"�	����u�֪,�/tM��楱����b��1ig!NN�0�z��(��,�.�
�ɺ?�#	*]]�iI9�o«IX0F�MSt�
���q���̰�!@EZ�����q9+t�}x��7�ֻ\1^O�Z�_v(��ƍ2���l���$PC�A�a��!/^�פ+��6��+�3�ET��;�jmT�#?�����&*rB�WD�{͘6��q����1ig!Ir��͕� h�ҩ�ݑ���&�d�+��\��F�̃��H��}Dq�f���Ě���ž_�F�(*�O�qs�۶��Z���>e�p�c)C�+�B-�DP����p��ݚ�Н�(@X~�H:5irAz.ln��뾦�!�`�(i3�5ߧE4���ݚ�Н����P� ^g�)�.�{�Y�Y�1!�`�(i3 �bVfj��h�c,.J���N���!�`�(i3�(R\֎u����>^17��"��ӌ�r���%>�rGO�D mWN;�jmT�#?�����&*rB�WD�{͘6��q����1ig!=�9E��@�� h�ҩ�ݑ���&�d�+��\��F�̃��H��}Dq�f���Ě���ž_�F�(*�O�q+y���,R�xB�<<۲��>e�p�c)C�+�B-�D(���27:����Kf��w�n9�gg��4p��o�+�B-�DP����p��ݚ�Н�(@X~�H:5irAz.ln��뾦�!�`�(i3�5ߧE4��!�`�(i3 �bVfj��h�c,.J�AԢ�a\�%o�P��(� ��0� 1tSjv���+�t2��\1^O�Z�_v(���?D�8��HN��R��F F�E̠ʁ���Mյ$��Q��@&U�)j�S���̰�!@EZ�����q9+t�}�ݚ�Н��(R\֎u�k�n�=���b+}y[�mJ�0�6�fĉ>99��|��3�W?�;�끶���A�����7�Y�Qqw�}�t����M~V��	��y ��f"�N#~8"�Z�<O�e�TL��c>d�xὕ?�5�e���Jm�W�)���䯐<!�̚��Ws� QӀ)&l�d�c�<���Lɓ6�C!c�"�ډ�.�n|����O�\0��6?�d���&�[��N�黬b��MF�̃��H��*k�Ҟv.�
�ɺ�)_�32����r����!�`�(i3���D4FF�v�����\1^O�Z�_v(��ڥ����Ⱦ��V8zA�o��<���� ��V��G��<��
ڰb��Ƽ��r����!�`�(i3���D4FF*���́;��|B���o1����-��uv=_j.;����e�
�J�s���:�H�+yx��Q��z�,�ML��e)����k�|��	>>E���O�m���Sc~��F�ET��ŢquA0�e]'\gWg��	�Z�kfcj��r���(&�L��'ž1�|��P�:k& ��-����N
����#�+#��]!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^��;��L�ז�1�, �y�`��vN1tSjv�7�wtMMiS���l�
���|e"���F��O�}�	76�&�� Ӗ�t$�)�vx.F<!W���2{��7��
����x���W�
�am�7#1=��*�����z��](g���М��^���'ƃ�3�Y�U��֯r~�p��8�5я����h�&�a�l����А����H�v�i�W��ɇ���J�4�KXh��`��1���~!�`�(i3��ӷ�*[D��:�%ЇD���Ѧ��*f1�.��N����k$ !�`�(i3��&j	Q�w�T� �f&���#��uގF1he��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc!N�'�y�G