��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���GK�趹���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�LZ*IV��ӓ�������]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R����h�K�5���� ��1�:�Ω�=A���>�LZ*IV��ӓ�������]P*m����)O��Ξ4�"�\�� ���K�O�{��?f���ʈj��U�sqc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c,� � U�rN�3��m-�@xI+r�� 0�D�A�f�mX��VNF��SK��1�����o�T�Y��6�J�|(���N�uD��N�uD��N�uD�_���TF�N�uD�_���TF_���TFWTd�'\q!�`�(i3��u�!�`�(i3��u�!�`�(i3��u�4�a�
�Ǜ��`$T)�	�
޼��	�
޼���G���s��z�*	.��G���s��4A��a_8|��K{l�+ׇӭ��!�`�(i3Jy�|�!�`�(i3!�`�(i3!�`�(i3,��L���!�`�(i3 ���M��mu�)L�!�`�(i3!�`�(i3�+���4ׇӭ��!�`�(i3!�`�(i3!�`�(i3g��A*	��!�`�(i3!�`�(i3!�`�(i3�+���4�WOtl��M!�nz��m��+��jTʱ�8F0_H��w�Sjs���N<��;���u��w)�S��X3����~篟|��
O�:��t����;r8�:r&@1�+Q�<��d���L!ۤՀ/Q9*سBK-����s~�j1���u��w)�S��X3�����@��."�;r|@�b�؃��em�J�Й�m��JNu���]�ߏ��P�umSe��S�2�:,�nr#�9l$�/P��pO�c�c�ENk�lAc>b�G��8̀@��k.�"SӠ�|&��c���m�Rܙ#l�%q�M�4�}�����r�N�Þ��t�U�PD@��k.͇�@�L�v���0�Rc=���T�1�\�^6uk��~1f��t�jPP�
� �AH����e��'�Wا[~�l]ǜ�����] ��F@�4%���D�Pfc����2P����/�"��< ���X�M+��tc��P9P��`�.�D���J7"9�x@�vD�t��⫓���RL�a))�kc�߇Bg�3���M Ce=6�([a�EF��7C��Hwɶ R�p��4�s4�o�qR��p������M<D�7�s)	w�N\`�a���!4d���-sk �0%̄sb�� bL�k>F�泂�0�V�@���RL�a)'r�Ӟh� mߍu�M9ts{z>�z�՝�ydѦ�7C��H!�������0�"���L�M�=o����"���	x]�
].~�Z�c�J�M=.��Ȁ�3���8�:r&@9����D��rG�K����B�6�*����	B�B��kQ����X���f+���J�J]�j�j�Ͼi0�?�"���D��(�1C`��^�1����2��BX��w-�����:��*����	�v`)��D��竺q�	r�O��C��0��?,*���S�K�?g�W"��!�1\Z��uDp�7C��H�z�/�E���d/^���,��:N�F&�Lki�Ijg��T��`e�:�$�i��Ahh](鞎�cX<����!�p�Ԉ��o�m�<H@���u�7X�K0o�6=� ������J c��(�U����	x]�m�Je{q��N��(
{��DIU�J���<���&}Xa���������dG�b�{����V���	x]���Ec��$7��Mv�9��!��|�����dC<8�:r&@L���Qep��p�R��$���wT��xݣL����RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QLi/-�#�v-~x��䂁!�o��c��(r���U����+rb�SO,F=d9�[l�&��q�©���H��JnXe�+�Uz�QLi/-�#�^ �Y�)��H*�m���b��y�.V&��B֥�(����5���I�zI.��1��bL�Y�͋�<Ct�z&��ÃlO ܅d^�R@Κ�2���ei"�,�>E����\�vňu�,�s�^�R@Κ�2�l~�Uf���}��\�v�T?�7G|`�UxHj,��|��	�"�,�>E����\�vňu�,�s���2��̪U��֜��3"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3JHn��z�_c)���8���bg�1�Z���=�������b9����,����d���z���ߘ�)�I��<
DN�l0��F��j�q	k���A���������]c���H������i�=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3���D	��U�l>o��|�,+$\�M��wF4��0[����	��N�Ae�#����ꀍ!�`�(i3c��Et��q���U����?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-�|�)՜�4!�`�(i3v�ј�"��Z鎬����(��eظ�_--���g&e�l�����-��%Mm�jp=�>��o�
�v�ξ������ei]��fM?R�^Ƒ����"X��[��Q[R�7W����GS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l����G<�e��
T�v��1���6��	���`y����ꢤ�OgZ)[���F�����E��@IE�U��n�-�6��
�jW��D���M���R'),��`��{|*�"��i�_:���5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f�ja1�n�[�c�/�O��?�;��XC�g����<ë��r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+��jTʱ�8F0_H��w�Sjs���-;���:��#I�90gA�I�y�?ܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'��!�a��5�%]���a(􆿳��?ƾ�؀qjZ��H@H�֦g�㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���o���ia���lC��U�T�\ ��y�.�`L⯆�'��wb�*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85��p#�j\1�Z���=�"j���b7|#9���b!��u��<��>��hs5e�U!K��tf��
_�n�@/%{�;����f�kN�ı&l����[}�@��L}�
�?��u��g��L`��Lל��[��Q�՝�i�(�S��]Q�I����踫g(�r� k�|6�8-+��B�G����n9��
����Ş��'^��\|YX�<I@1�ؠ&���Z02�	L�E����Y�7#�xI�_II� �*��H��,Q���36�`��������8�QuXu�[pUI��'��d�uY��dzw⭏l�u��s$y�<5������U��֜��3��P=@��������$��Xo�-��8�%���ތ�1�"5� �S��eP�Y�7#�xIG�2ƨ�ܠ����\��0���1�(�����@^7&ģM��`�z��GZ>.�0�XpɽP��a�x��d�uY�ا�W��_�ړ8���/�I����"��T:���V������?�7�>l�r�z*���Be�2l��4��a��se�ξ������ei4����/��)}���/��r��H��g��m������H���	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8�	�A��ԡe���b�kvo�Apw��0���1���@c
�YqJH��[q�t��c_����+�˂߮<uȧh}�ulj��^̽1�� k�|6�8�Qe�`�=`<�Fk R- j�i�+-�6��.��L�L;Л��|#9�����w��l�oP��a�I�;��0���}����g������h^:�髊}�B�]��871��B�D�F v��[6"����|!�^����N>�4�
��i��,�/����~9��4�듴,`Y�{'%s4���"�wq�0B��f'?	G݈�����a�"Z鎬�������(��`UNP� ��b�FP&���P��'���Xw�j�7���1�L�+��8���/��8&���I��I�Cp�GEE�ޱ� p-�a &r|�t�iiTqm5|X������[ Ӄ2�R����������t�'jf�|sb�d"L�Ɯd� (�f퀔����`0�S�����N�|�("0�i��$��lq�0�+��J@�h�����XX���Ě�����������E@=�>�V�Re��Q�8���/�T���Pk�7�癆cg���K�Ou�0��uϊ���v�қp �u��r��7�%M��4f�x #^�9n��,�J��/3o�U�r*A&-�Ri֭�h��O��@�D%����6Q���,G�_baHN��R���מu��� �H�0��
1���~��=�g���>��i)�'a>-#�}�7��[��(���y��j��kj�����N�/��kOT���W0�]��e|)0�٣ԩ|���}�	76�&��A0ok��6�������ݸ���TT7���1����#M&�4�q�Xx�=�6%j_�zJe��0��-&�6��_���9�j�u���G5�O�%E#P�≯
�Ϗ�i7N�_�z*K�/��=��K�9T��,�����Z��!�`�(i3'G�+R���o��_�Rv�䩲$���dS@Ɵ�o��6}���(&�L�;�jmT�#bs��2[�a��o���H�RtV�^�2��}�������Ə��.A`��x��nF���<�W�.�P�	��
�Q�}!�`�(i3mj�B��Vh�EtC�<�b_X�XV�b�z'hۉ)��d�7�q�!�`�(i3)�{6�U���Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#!�`�(i3܌;���'����u��r��!�`�(i3��TBd��pS�*;q܆QCj�4Z�_--���gz���M�~}!�`�(i3�G�dE�h�����?uA|�d���u��g��L�}M�9s��!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rG߸��S�Ȍ����PJfĉ>99��;��|B	���>o��.�g3ZE��g�Hb�? tB&�kM�����y48{���@2P�)�#�Xgjn3ԏ�W+��W���TBd��pS�*;q�v{��lw	�,Bp��S���.J7h��r��H�Cw�Hm��mj�B��Vφ�?'�Q����,�ǰ��i��W�o`�k�������.ʀ8�t�|2;$�JأͽgF"?�Q��ǺΕ�f�f3'_��s�֙Ш��"x���������o��_�Rv�䩲$���dS@Ɵ�od=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^��4-�b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu��� ߛ��usȸ�"rR��U��3i�z6��s�u��p��V�M'��w]Pi�#��R!�`�(i3=��,���H̷_��yC��S8�����ZK����t����>3���w�@V-���,W������0�� 7�J�[|�m�ߕ��[���#�!�`�(i3�Y�m�k?j!�`�(i3�/�cLbŪ�����:Y�{'%s��$��S���b�Bϱ��<��>��h�EtC�<�+������L�*dgN;�r��H�?X���V4&v��؄aX�
�:qEp�;�P�t�5!�`�(i37�A��\R��c���鿡�t����>3���w�@V-���,W������0�� 7�J�[|�m�ߕ��:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6���@P?�(w�R���y�sL]~цߒ�a`p�Y�u7B�k"-�i7N�_�Ar��� ����Dɵ�p�AJ�e�$��8y�Ɋ����Z��d�G}%��Ď��J��QCT�"�x9�¿Y�����ϪE�smy^� 3�hD�p~z�r,wK��-��}��d���!i�SENan&�������%q�>��8�>r&���c
� ��;��|B���r��������o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!q��V���<	s/.�Ss�g��+˘\5���jmY�VS���g�n�{�6�e
��>�i�g��+˘\5���jmY��X"e_�4�{�6�em�;���HN��R��?�d���&��Ebu��SENan&�\�0Iѓ�1M� Ѯ&U��8�>r&��U������yf��>5�O�%E#PZt%��m&<�P8��PS~�Dn��i�Q׭n�L���/=9j���)��Q��\@
��:�)�<�����⪂!t-�u	D�&���A3�Q��\@
����G3҇
��'T���+`��W#s�2t�N�/�ڃ����<N߼�K�iN�� ��Tv-_�0!>���@]��}Dq�f�����,�ǰE��C$�����B���'�綅������>vD���&l����$�<�F�q;��|B���r��������o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!q��V���<	s/����AIe��0�U+�qbp@����%>�rG6j�"Hs��}�R�s���Z/���Bj���!�9ה;�Q��ǺΕod'ٙ� �z�:Y���J��:����SƏw0��C�ݥc&���XO)�Q>�W��*(��3H��ieL���1��#��{�6�em�;���Zt%��m&<�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��pw�R���y��0�J���B:�cV��	��yv�ʯʗYo��g��N�1��#�s��e�i��ƫg�T�k�Y���;��|B���r�������`3�Jg'X�~bw��U��)���Y;e�iK!���d.[�����:Fa�7��-Ukc��R2�e��b�uz۴k1��˪���l��A(�c���_G��Hb� h�ҩ�SƏw0��C�ݥc&���XO)�Q�{_8�Y��=�}�Vݨ��}Dq�f�FkH��۟�z��n� ���?R �K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��=�O�-v�*_�mS8<�n�ݚ�Н��H����Q�R���F�(|��8����ei�B� �b��!�`�(i3SƏw0��C�ݥc&���XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���!�`�(i3FkH��۟�z��n� ���?R �����⪂!t-�u	D�&F�WAM�Q��\@
��:�)�<�����⪂!t-�u	D�&6���G1�Q��\@
����G3҇
!�`�(i3�̢k���:�ct�0��3��O	�T/ k�|6�878�^9u��r��!�`�(i3����o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!�`�(i3��hY-N�g3�)��c�{I���,'�*;���#�b�>{Z����6��.��Lj�)6)-
!�`�(i3>��iC���D����_ �Q��ǺΕod'ٙ� �~��<e�3�ݚ�Н���'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3Zt%��m&<�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��p
�:qEp'{w#/ B!�`�(i3����o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ��:5A��p!�`�(i3��hY-N�g3�)��b_X�XV�b�z'hۉ)��d�7�q�!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Fr��j~�8�r\���1 ��b�i3�I��)���W�w��fD^����+���F�}қ~�C탤ϻ�U��)���Y;e�iKI/B޾PԐ#��go`iI9�o��|#HK��A(�c���_G��Hb� h�ҩ�!q��V��w:��<����nF���<�W�.�P�	��
�Q�}�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��
�t��T&���LQ�/81tSjv���'T���+�E���v��g����`��W#s�m4V2�@�P8��PS~��Q���N�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jr��*�tB+p�^(w�R���y"O���%jm
�����"�7�\�`,9�H�W��`�z6/������,���eFz�qb	��G��W+��W��.W��&k@C�Ɨ0z�cUL��Zi+�E��ĵ�%�'�֝�p6j�"Hsۍ=Z�&�Jƨ�Jt̫j(&
M�K;��%YM�	�v�3� k�|6�8��:�EB�Z5�O�%E#P#L�
�am$��	��#�|����m�I7��-55x|���MM
��,=?�d���&�t�{#	�x��_--���g�QF.��v{��lw	�����?QZ���>��,H/������,�ǰ�������Z���zh�#L�
�am$�Z�^��h�@^4KT�v��1�5x|���MM
��,=?�d���&���=����t 7�J�[> a��M����DKY�������?QZ���>ś���k�����,�ǰ�������m2�
��E����,�ǰu!�OO��
}Z8/��RU��H��<�C�Ar��� ����Dɵ�p�AJ�e�$��8y�Ɋ����Z���F%�X��k��o������"O��_U)�<�&#R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0�`j3���Fm�b�vA`v@񴱝�P���Q�w�R���ykb>���pP�|x����.�g3Zdj�t��C���j��~(㷾�N���H݆�